module bht(
  input         clock,
  input         reset,
  input         io_valid,
  input  [31:0] io_pc,
  output        io_takenPre,
  output        io_ready,
  input         io_takenValid,
  input         io_takenMiss,
  input         io_exTakenPre,
  input  [31:0] io_takenPC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ghr; // @[bht.scala 51:22]
  reg [7:0] bht_0; // @[bht.scala 52:22]
  reg [7:0] bht_1; // @[bht.scala 52:22]
  reg [7:0] bht_2; // @[bht.scala 52:22]
  reg [7:0] bht_3; // @[bht.scala 52:22]
  reg [7:0] bht_4; // @[bht.scala 52:22]
  reg [7:0] bht_5; // @[bht.scala 52:22]
  reg [7:0] bht_6; // @[bht.scala 52:22]
  reg [7:0] bht_7; // @[bht.scala 52:22]
  reg [7:0] bht_8; // @[bht.scala 52:22]
  reg [7:0] bht_9; // @[bht.scala 52:22]
  reg [7:0] bht_10; // @[bht.scala 52:22]
  reg [7:0] bht_11; // @[bht.scala 52:22]
  reg [7:0] bht_12; // @[bht.scala 52:22]
  reg [7:0] bht_13; // @[bht.scala 52:22]
  reg [7:0] bht_14; // @[bht.scala 52:22]
  reg [7:0] bht_15; // @[bht.scala 52:22]
  reg [7:0] bht_16; // @[bht.scala 52:22]
  reg [7:0] bht_17; // @[bht.scala 52:22]
  reg [7:0] bht_18; // @[bht.scala 52:22]
  reg [7:0] bht_19; // @[bht.scala 52:22]
  reg [7:0] bht_20; // @[bht.scala 52:22]
  reg [7:0] bht_21; // @[bht.scala 52:22]
  reg [7:0] bht_22; // @[bht.scala 52:22]
  reg [7:0] bht_23; // @[bht.scala 52:22]
  reg [7:0] bht_24; // @[bht.scala 52:22]
  reg [7:0] bht_25; // @[bht.scala 52:22]
  reg [7:0] bht_26; // @[bht.scala 52:22]
  reg [7:0] bht_27; // @[bht.scala 52:22]
  reg [7:0] bht_28; // @[bht.scala 52:22]
  reg [7:0] bht_29; // @[bht.scala 52:22]
  reg [7:0] bht_30; // @[bht.scala 52:22]
  reg [7:0] bht_31; // @[bht.scala 52:22]
  reg [7:0] bht_32; // @[bht.scala 52:22]
  reg [7:0] bht_33; // @[bht.scala 52:22]
  reg [7:0] bht_34; // @[bht.scala 52:22]
  reg [7:0] bht_35; // @[bht.scala 52:22]
  reg [7:0] bht_36; // @[bht.scala 52:22]
  reg [7:0] bht_37; // @[bht.scala 52:22]
  reg [7:0] bht_38; // @[bht.scala 52:22]
  reg [7:0] bht_39; // @[bht.scala 52:22]
  reg [7:0] bht_40; // @[bht.scala 52:22]
  reg [7:0] bht_41; // @[bht.scala 52:22]
  reg [7:0] bht_42; // @[bht.scala 52:22]
  reg [7:0] bht_43; // @[bht.scala 52:22]
  reg [7:0] bht_44; // @[bht.scala 52:22]
  reg [7:0] bht_45; // @[bht.scala 52:22]
  reg [7:0] bht_46; // @[bht.scala 52:22]
  reg [7:0] bht_47; // @[bht.scala 52:22]
  reg [7:0] bht_48; // @[bht.scala 52:22]
  reg [7:0] bht_49; // @[bht.scala 52:22]
  reg [7:0] bht_50; // @[bht.scala 52:22]
  reg [7:0] bht_51; // @[bht.scala 52:22]
  reg [7:0] bht_52; // @[bht.scala 52:22]
  reg [7:0] bht_53; // @[bht.scala 52:22]
  reg [7:0] bht_54; // @[bht.scala 52:22]
  reg [7:0] bht_55; // @[bht.scala 52:22]
  reg [7:0] bht_56; // @[bht.scala 52:22]
  reg [7:0] bht_57; // @[bht.scala 52:22]
  reg [7:0] bht_58; // @[bht.scala 52:22]
  reg [7:0] bht_59; // @[bht.scala 52:22]
  reg [7:0] bht_60; // @[bht.scala 52:22]
  reg [7:0] bht_61; // @[bht.scala 52:22]
  reg [7:0] bht_62; // @[bht.scala 52:22]
  reg [7:0] bht_63; // @[bht.scala 52:22]
  reg [1:0] pht_0_0; // @[bht.scala 53:22]
  reg [1:0] pht_0_1; // @[bht.scala 53:22]
  reg [1:0] pht_0_2; // @[bht.scala 53:22]
  reg [1:0] pht_0_3; // @[bht.scala 53:22]
  reg [1:0] pht_0_4; // @[bht.scala 53:22]
  reg [1:0] pht_0_5; // @[bht.scala 53:22]
  reg [1:0] pht_0_6; // @[bht.scala 53:22]
  reg [1:0] pht_0_7; // @[bht.scala 53:22]
  reg [1:0] pht_0_8; // @[bht.scala 53:22]
  reg [1:0] pht_0_9; // @[bht.scala 53:22]
  reg [1:0] pht_0_10; // @[bht.scala 53:22]
  reg [1:0] pht_0_11; // @[bht.scala 53:22]
  reg [1:0] pht_0_12; // @[bht.scala 53:22]
  reg [1:0] pht_0_13; // @[bht.scala 53:22]
  reg [1:0] pht_0_14; // @[bht.scala 53:22]
  reg [1:0] pht_0_15; // @[bht.scala 53:22]
  reg [1:0] pht_0_16; // @[bht.scala 53:22]
  reg [1:0] pht_0_17; // @[bht.scala 53:22]
  reg [1:0] pht_0_18; // @[bht.scala 53:22]
  reg [1:0] pht_0_19; // @[bht.scala 53:22]
  reg [1:0] pht_0_20; // @[bht.scala 53:22]
  reg [1:0] pht_0_21; // @[bht.scala 53:22]
  reg [1:0] pht_0_22; // @[bht.scala 53:22]
  reg [1:0] pht_0_23; // @[bht.scala 53:22]
  reg [1:0] pht_0_24; // @[bht.scala 53:22]
  reg [1:0] pht_0_25; // @[bht.scala 53:22]
  reg [1:0] pht_0_26; // @[bht.scala 53:22]
  reg [1:0] pht_0_27; // @[bht.scala 53:22]
  reg [1:0] pht_0_28; // @[bht.scala 53:22]
  reg [1:0] pht_0_29; // @[bht.scala 53:22]
  reg [1:0] pht_0_30; // @[bht.scala 53:22]
  reg [1:0] pht_0_31; // @[bht.scala 53:22]
  reg [1:0] pht_0_32; // @[bht.scala 53:22]
  reg [1:0] pht_0_33; // @[bht.scala 53:22]
  reg [1:0] pht_0_34; // @[bht.scala 53:22]
  reg [1:0] pht_0_35; // @[bht.scala 53:22]
  reg [1:0] pht_0_36; // @[bht.scala 53:22]
  reg [1:0] pht_0_37; // @[bht.scala 53:22]
  reg [1:0] pht_0_38; // @[bht.scala 53:22]
  reg [1:0] pht_0_39; // @[bht.scala 53:22]
  reg [1:0] pht_0_40; // @[bht.scala 53:22]
  reg [1:0] pht_0_41; // @[bht.scala 53:22]
  reg [1:0] pht_0_42; // @[bht.scala 53:22]
  reg [1:0] pht_0_43; // @[bht.scala 53:22]
  reg [1:0] pht_0_44; // @[bht.scala 53:22]
  reg [1:0] pht_0_45; // @[bht.scala 53:22]
  reg [1:0] pht_0_46; // @[bht.scala 53:22]
  reg [1:0] pht_0_47; // @[bht.scala 53:22]
  reg [1:0] pht_0_48; // @[bht.scala 53:22]
  reg [1:0] pht_0_49; // @[bht.scala 53:22]
  reg [1:0] pht_0_50; // @[bht.scala 53:22]
  reg [1:0] pht_0_51; // @[bht.scala 53:22]
  reg [1:0] pht_0_52; // @[bht.scala 53:22]
  reg [1:0] pht_0_53; // @[bht.scala 53:22]
  reg [1:0] pht_0_54; // @[bht.scala 53:22]
  reg [1:0] pht_0_55; // @[bht.scala 53:22]
  reg [1:0] pht_0_56; // @[bht.scala 53:22]
  reg [1:0] pht_0_57; // @[bht.scala 53:22]
  reg [1:0] pht_0_58; // @[bht.scala 53:22]
  reg [1:0] pht_0_59; // @[bht.scala 53:22]
  reg [1:0] pht_0_60; // @[bht.scala 53:22]
  reg [1:0] pht_0_61; // @[bht.scala 53:22]
  reg [1:0] pht_0_62; // @[bht.scala 53:22]
  reg [1:0] pht_0_63; // @[bht.scala 53:22]
  reg [1:0] pht_0_64; // @[bht.scala 53:22]
  reg [1:0] pht_0_65; // @[bht.scala 53:22]
  reg [1:0] pht_0_66; // @[bht.scala 53:22]
  reg [1:0] pht_0_67; // @[bht.scala 53:22]
  reg [1:0] pht_0_68; // @[bht.scala 53:22]
  reg [1:0] pht_0_69; // @[bht.scala 53:22]
  reg [1:0] pht_0_70; // @[bht.scala 53:22]
  reg [1:0] pht_0_71; // @[bht.scala 53:22]
  reg [1:0] pht_0_72; // @[bht.scala 53:22]
  reg [1:0] pht_0_73; // @[bht.scala 53:22]
  reg [1:0] pht_0_74; // @[bht.scala 53:22]
  reg [1:0] pht_0_75; // @[bht.scala 53:22]
  reg [1:0] pht_0_76; // @[bht.scala 53:22]
  reg [1:0] pht_0_77; // @[bht.scala 53:22]
  reg [1:0] pht_0_78; // @[bht.scala 53:22]
  reg [1:0] pht_0_79; // @[bht.scala 53:22]
  reg [1:0] pht_0_80; // @[bht.scala 53:22]
  reg [1:0] pht_0_81; // @[bht.scala 53:22]
  reg [1:0] pht_0_82; // @[bht.scala 53:22]
  reg [1:0] pht_0_83; // @[bht.scala 53:22]
  reg [1:0] pht_0_84; // @[bht.scala 53:22]
  reg [1:0] pht_0_85; // @[bht.scala 53:22]
  reg [1:0] pht_0_86; // @[bht.scala 53:22]
  reg [1:0] pht_0_87; // @[bht.scala 53:22]
  reg [1:0] pht_0_88; // @[bht.scala 53:22]
  reg [1:0] pht_0_89; // @[bht.scala 53:22]
  reg [1:0] pht_0_90; // @[bht.scala 53:22]
  reg [1:0] pht_0_91; // @[bht.scala 53:22]
  reg [1:0] pht_0_92; // @[bht.scala 53:22]
  reg [1:0] pht_0_93; // @[bht.scala 53:22]
  reg [1:0] pht_0_94; // @[bht.scala 53:22]
  reg [1:0] pht_0_95; // @[bht.scala 53:22]
  reg [1:0] pht_0_96; // @[bht.scala 53:22]
  reg [1:0] pht_0_97; // @[bht.scala 53:22]
  reg [1:0] pht_0_98; // @[bht.scala 53:22]
  reg [1:0] pht_0_99; // @[bht.scala 53:22]
  reg [1:0] pht_0_100; // @[bht.scala 53:22]
  reg [1:0] pht_0_101; // @[bht.scala 53:22]
  reg [1:0] pht_0_102; // @[bht.scala 53:22]
  reg [1:0] pht_0_103; // @[bht.scala 53:22]
  reg [1:0] pht_0_104; // @[bht.scala 53:22]
  reg [1:0] pht_0_105; // @[bht.scala 53:22]
  reg [1:0] pht_0_106; // @[bht.scala 53:22]
  reg [1:0] pht_0_107; // @[bht.scala 53:22]
  reg [1:0] pht_0_108; // @[bht.scala 53:22]
  reg [1:0] pht_0_109; // @[bht.scala 53:22]
  reg [1:0] pht_0_110; // @[bht.scala 53:22]
  reg [1:0] pht_0_111; // @[bht.scala 53:22]
  reg [1:0] pht_0_112; // @[bht.scala 53:22]
  reg [1:0] pht_0_113; // @[bht.scala 53:22]
  reg [1:0] pht_0_114; // @[bht.scala 53:22]
  reg [1:0] pht_0_115; // @[bht.scala 53:22]
  reg [1:0] pht_0_116; // @[bht.scala 53:22]
  reg [1:0] pht_0_117; // @[bht.scala 53:22]
  reg [1:0] pht_0_118; // @[bht.scala 53:22]
  reg [1:0] pht_0_119; // @[bht.scala 53:22]
  reg [1:0] pht_0_120; // @[bht.scala 53:22]
  reg [1:0] pht_0_121; // @[bht.scala 53:22]
  reg [1:0] pht_0_122; // @[bht.scala 53:22]
  reg [1:0] pht_0_123; // @[bht.scala 53:22]
  reg [1:0] pht_0_124; // @[bht.scala 53:22]
  reg [1:0] pht_0_125; // @[bht.scala 53:22]
  reg [1:0] pht_0_126; // @[bht.scala 53:22]
  reg [1:0] pht_0_127; // @[bht.scala 53:22]
  reg [1:0] pht_0_128; // @[bht.scala 53:22]
  reg [1:0] pht_0_129; // @[bht.scala 53:22]
  reg [1:0] pht_0_130; // @[bht.scala 53:22]
  reg [1:0] pht_0_131; // @[bht.scala 53:22]
  reg [1:0] pht_0_132; // @[bht.scala 53:22]
  reg [1:0] pht_0_133; // @[bht.scala 53:22]
  reg [1:0] pht_0_134; // @[bht.scala 53:22]
  reg [1:0] pht_0_135; // @[bht.scala 53:22]
  reg [1:0] pht_0_136; // @[bht.scala 53:22]
  reg [1:0] pht_0_137; // @[bht.scala 53:22]
  reg [1:0] pht_0_138; // @[bht.scala 53:22]
  reg [1:0] pht_0_139; // @[bht.scala 53:22]
  reg [1:0] pht_0_140; // @[bht.scala 53:22]
  reg [1:0] pht_0_141; // @[bht.scala 53:22]
  reg [1:0] pht_0_142; // @[bht.scala 53:22]
  reg [1:0] pht_0_143; // @[bht.scala 53:22]
  reg [1:0] pht_0_144; // @[bht.scala 53:22]
  reg [1:0] pht_0_145; // @[bht.scala 53:22]
  reg [1:0] pht_0_146; // @[bht.scala 53:22]
  reg [1:0] pht_0_147; // @[bht.scala 53:22]
  reg [1:0] pht_0_148; // @[bht.scala 53:22]
  reg [1:0] pht_0_149; // @[bht.scala 53:22]
  reg [1:0] pht_0_150; // @[bht.scala 53:22]
  reg [1:0] pht_0_151; // @[bht.scala 53:22]
  reg [1:0] pht_0_152; // @[bht.scala 53:22]
  reg [1:0] pht_0_153; // @[bht.scala 53:22]
  reg [1:0] pht_0_154; // @[bht.scala 53:22]
  reg [1:0] pht_0_155; // @[bht.scala 53:22]
  reg [1:0] pht_0_156; // @[bht.scala 53:22]
  reg [1:0] pht_0_157; // @[bht.scala 53:22]
  reg [1:0] pht_0_158; // @[bht.scala 53:22]
  reg [1:0] pht_0_159; // @[bht.scala 53:22]
  reg [1:0] pht_0_160; // @[bht.scala 53:22]
  reg [1:0] pht_0_161; // @[bht.scala 53:22]
  reg [1:0] pht_0_162; // @[bht.scala 53:22]
  reg [1:0] pht_0_163; // @[bht.scala 53:22]
  reg [1:0] pht_0_164; // @[bht.scala 53:22]
  reg [1:0] pht_0_165; // @[bht.scala 53:22]
  reg [1:0] pht_0_166; // @[bht.scala 53:22]
  reg [1:0] pht_0_167; // @[bht.scala 53:22]
  reg [1:0] pht_0_168; // @[bht.scala 53:22]
  reg [1:0] pht_0_169; // @[bht.scala 53:22]
  reg [1:0] pht_0_170; // @[bht.scala 53:22]
  reg [1:0] pht_0_171; // @[bht.scala 53:22]
  reg [1:0] pht_0_172; // @[bht.scala 53:22]
  reg [1:0] pht_0_173; // @[bht.scala 53:22]
  reg [1:0] pht_0_174; // @[bht.scala 53:22]
  reg [1:0] pht_0_175; // @[bht.scala 53:22]
  reg [1:0] pht_0_176; // @[bht.scala 53:22]
  reg [1:0] pht_0_177; // @[bht.scala 53:22]
  reg [1:0] pht_0_178; // @[bht.scala 53:22]
  reg [1:0] pht_0_179; // @[bht.scala 53:22]
  reg [1:0] pht_0_180; // @[bht.scala 53:22]
  reg [1:0] pht_0_181; // @[bht.scala 53:22]
  reg [1:0] pht_0_182; // @[bht.scala 53:22]
  reg [1:0] pht_0_183; // @[bht.scala 53:22]
  reg [1:0] pht_0_184; // @[bht.scala 53:22]
  reg [1:0] pht_0_185; // @[bht.scala 53:22]
  reg [1:0] pht_0_186; // @[bht.scala 53:22]
  reg [1:0] pht_0_187; // @[bht.scala 53:22]
  reg [1:0] pht_0_188; // @[bht.scala 53:22]
  reg [1:0] pht_0_189; // @[bht.scala 53:22]
  reg [1:0] pht_0_190; // @[bht.scala 53:22]
  reg [1:0] pht_0_191; // @[bht.scala 53:22]
  reg [1:0] pht_0_192; // @[bht.scala 53:22]
  reg [1:0] pht_0_193; // @[bht.scala 53:22]
  reg [1:0] pht_0_194; // @[bht.scala 53:22]
  reg [1:0] pht_0_195; // @[bht.scala 53:22]
  reg [1:0] pht_0_196; // @[bht.scala 53:22]
  reg [1:0] pht_0_197; // @[bht.scala 53:22]
  reg [1:0] pht_0_198; // @[bht.scala 53:22]
  reg [1:0] pht_0_199; // @[bht.scala 53:22]
  reg [1:0] pht_0_200; // @[bht.scala 53:22]
  reg [1:0] pht_0_201; // @[bht.scala 53:22]
  reg [1:0] pht_0_202; // @[bht.scala 53:22]
  reg [1:0] pht_0_203; // @[bht.scala 53:22]
  reg [1:0] pht_0_204; // @[bht.scala 53:22]
  reg [1:0] pht_0_205; // @[bht.scala 53:22]
  reg [1:0] pht_0_206; // @[bht.scala 53:22]
  reg [1:0] pht_0_207; // @[bht.scala 53:22]
  reg [1:0] pht_0_208; // @[bht.scala 53:22]
  reg [1:0] pht_0_209; // @[bht.scala 53:22]
  reg [1:0] pht_0_210; // @[bht.scala 53:22]
  reg [1:0] pht_0_211; // @[bht.scala 53:22]
  reg [1:0] pht_0_212; // @[bht.scala 53:22]
  reg [1:0] pht_0_213; // @[bht.scala 53:22]
  reg [1:0] pht_0_214; // @[bht.scala 53:22]
  reg [1:0] pht_0_215; // @[bht.scala 53:22]
  reg [1:0] pht_0_216; // @[bht.scala 53:22]
  reg [1:0] pht_0_217; // @[bht.scala 53:22]
  reg [1:0] pht_0_218; // @[bht.scala 53:22]
  reg [1:0] pht_0_219; // @[bht.scala 53:22]
  reg [1:0] pht_0_220; // @[bht.scala 53:22]
  reg [1:0] pht_0_221; // @[bht.scala 53:22]
  reg [1:0] pht_0_222; // @[bht.scala 53:22]
  reg [1:0] pht_0_223; // @[bht.scala 53:22]
  reg [1:0] pht_0_224; // @[bht.scala 53:22]
  reg [1:0] pht_0_225; // @[bht.scala 53:22]
  reg [1:0] pht_0_226; // @[bht.scala 53:22]
  reg [1:0] pht_0_227; // @[bht.scala 53:22]
  reg [1:0] pht_0_228; // @[bht.scala 53:22]
  reg [1:0] pht_0_229; // @[bht.scala 53:22]
  reg [1:0] pht_0_230; // @[bht.scala 53:22]
  reg [1:0] pht_0_231; // @[bht.scala 53:22]
  reg [1:0] pht_0_232; // @[bht.scala 53:22]
  reg [1:0] pht_0_233; // @[bht.scala 53:22]
  reg [1:0] pht_0_234; // @[bht.scala 53:22]
  reg [1:0] pht_0_235; // @[bht.scala 53:22]
  reg [1:0] pht_0_236; // @[bht.scala 53:22]
  reg [1:0] pht_0_237; // @[bht.scala 53:22]
  reg [1:0] pht_0_238; // @[bht.scala 53:22]
  reg [1:0] pht_0_239; // @[bht.scala 53:22]
  reg [1:0] pht_0_240; // @[bht.scala 53:22]
  reg [1:0] pht_0_241; // @[bht.scala 53:22]
  reg [1:0] pht_0_242; // @[bht.scala 53:22]
  reg [1:0] pht_0_243; // @[bht.scala 53:22]
  reg [1:0] pht_0_244; // @[bht.scala 53:22]
  reg [1:0] pht_0_245; // @[bht.scala 53:22]
  reg [1:0] pht_0_246; // @[bht.scala 53:22]
  reg [1:0] pht_0_247; // @[bht.scala 53:22]
  reg [1:0] pht_0_248; // @[bht.scala 53:22]
  reg [1:0] pht_0_249; // @[bht.scala 53:22]
  reg [1:0] pht_0_250; // @[bht.scala 53:22]
  reg [1:0] pht_0_251; // @[bht.scala 53:22]
  reg [1:0] pht_0_252; // @[bht.scala 53:22]
  reg [1:0] pht_0_253; // @[bht.scala 53:22]
  reg [1:0] pht_0_254; // @[bht.scala 53:22]
  reg [1:0] pht_0_255; // @[bht.scala 53:22]
  reg [1:0] pht_1_0; // @[bht.scala 53:22]
  reg [1:0] pht_1_1; // @[bht.scala 53:22]
  reg [1:0] pht_1_2; // @[bht.scala 53:22]
  reg [1:0] pht_1_3; // @[bht.scala 53:22]
  reg [1:0] pht_1_4; // @[bht.scala 53:22]
  reg [1:0] pht_1_5; // @[bht.scala 53:22]
  reg [1:0] pht_1_6; // @[bht.scala 53:22]
  reg [1:0] pht_1_7; // @[bht.scala 53:22]
  reg [1:0] pht_1_8; // @[bht.scala 53:22]
  reg [1:0] pht_1_9; // @[bht.scala 53:22]
  reg [1:0] pht_1_10; // @[bht.scala 53:22]
  reg [1:0] pht_1_11; // @[bht.scala 53:22]
  reg [1:0] pht_1_12; // @[bht.scala 53:22]
  reg [1:0] pht_1_13; // @[bht.scala 53:22]
  reg [1:0] pht_1_14; // @[bht.scala 53:22]
  reg [1:0] pht_1_15; // @[bht.scala 53:22]
  reg [1:0] pht_1_16; // @[bht.scala 53:22]
  reg [1:0] pht_1_17; // @[bht.scala 53:22]
  reg [1:0] pht_1_18; // @[bht.scala 53:22]
  reg [1:0] pht_1_19; // @[bht.scala 53:22]
  reg [1:0] pht_1_20; // @[bht.scala 53:22]
  reg [1:0] pht_1_21; // @[bht.scala 53:22]
  reg [1:0] pht_1_22; // @[bht.scala 53:22]
  reg [1:0] pht_1_23; // @[bht.scala 53:22]
  reg [1:0] pht_1_24; // @[bht.scala 53:22]
  reg [1:0] pht_1_25; // @[bht.scala 53:22]
  reg [1:0] pht_1_26; // @[bht.scala 53:22]
  reg [1:0] pht_1_27; // @[bht.scala 53:22]
  reg [1:0] pht_1_28; // @[bht.scala 53:22]
  reg [1:0] pht_1_29; // @[bht.scala 53:22]
  reg [1:0] pht_1_30; // @[bht.scala 53:22]
  reg [1:0] pht_1_31; // @[bht.scala 53:22]
  reg [1:0] pht_1_32; // @[bht.scala 53:22]
  reg [1:0] pht_1_33; // @[bht.scala 53:22]
  reg [1:0] pht_1_34; // @[bht.scala 53:22]
  reg [1:0] pht_1_35; // @[bht.scala 53:22]
  reg [1:0] pht_1_36; // @[bht.scala 53:22]
  reg [1:0] pht_1_37; // @[bht.scala 53:22]
  reg [1:0] pht_1_38; // @[bht.scala 53:22]
  reg [1:0] pht_1_39; // @[bht.scala 53:22]
  reg [1:0] pht_1_40; // @[bht.scala 53:22]
  reg [1:0] pht_1_41; // @[bht.scala 53:22]
  reg [1:0] pht_1_42; // @[bht.scala 53:22]
  reg [1:0] pht_1_43; // @[bht.scala 53:22]
  reg [1:0] pht_1_44; // @[bht.scala 53:22]
  reg [1:0] pht_1_45; // @[bht.scala 53:22]
  reg [1:0] pht_1_46; // @[bht.scala 53:22]
  reg [1:0] pht_1_47; // @[bht.scala 53:22]
  reg [1:0] pht_1_48; // @[bht.scala 53:22]
  reg [1:0] pht_1_49; // @[bht.scala 53:22]
  reg [1:0] pht_1_50; // @[bht.scala 53:22]
  reg [1:0] pht_1_51; // @[bht.scala 53:22]
  reg [1:0] pht_1_52; // @[bht.scala 53:22]
  reg [1:0] pht_1_53; // @[bht.scala 53:22]
  reg [1:0] pht_1_54; // @[bht.scala 53:22]
  reg [1:0] pht_1_55; // @[bht.scala 53:22]
  reg [1:0] pht_1_56; // @[bht.scala 53:22]
  reg [1:0] pht_1_57; // @[bht.scala 53:22]
  reg [1:0] pht_1_58; // @[bht.scala 53:22]
  reg [1:0] pht_1_59; // @[bht.scala 53:22]
  reg [1:0] pht_1_60; // @[bht.scala 53:22]
  reg [1:0] pht_1_61; // @[bht.scala 53:22]
  reg [1:0] pht_1_62; // @[bht.scala 53:22]
  reg [1:0] pht_1_63; // @[bht.scala 53:22]
  reg [1:0] pht_1_64; // @[bht.scala 53:22]
  reg [1:0] pht_1_65; // @[bht.scala 53:22]
  reg [1:0] pht_1_66; // @[bht.scala 53:22]
  reg [1:0] pht_1_67; // @[bht.scala 53:22]
  reg [1:0] pht_1_68; // @[bht.scala 53:22]
  reg [1:0] pht_1_69; // @[bht.scala 53:22]
  reg [1:0] pht_1_70; // @[bht.scala 53:22]
  reg [1:0] pht_1_71; // @[bht.scala 53:22]
  reg [1:0] pht_1_72; // @[bht.scala 53:22]
  reg [1:0] pht_1_73; // @[bht.scala 53:22]
  reg [1:0] pht_1_74; // @[bht.scala 53:22]
  reg [1:0] pht_1_75; // @[bht.scala 53:22]
  reg [1:0] pht_1_76; // @[bht.scala 53:22]
  reg [1:0] pht_1_77; // @[bht.scala 53:22]
  reg [1:0] pht_1_78; // @[bht.scala 53:22]
  reg [1:0] pht_1_79; // @[bht.scala 53:22]
  reg [1:0] pht_1_80; // @[bht.scala 53:22]
  reg [1:0] pht_1_81; // @[bht.scala 53:22]
  reg [1:0] pht_1_82; // @[bht.scala 53:22]
  reg [1:0] pht_1_83; // @[bht.scala 53:22]
  reg [1:0] pht_1_84; // @[bht.scala 53:22]
  reg [1:0] pht_1_85; // @[bht.scala 53:22]
  reg [1:0] pht_1_86; // @[bht.scala 53:22]
  reg [1:0] pht_1_87; // @[bht.scala 53:22]
  reg [1:0] pht_1_88; // @[bht.scala 53:22]
  reg [1:0] pht_1_89; // @[bht.scala 53:22]
  reg [1:0] pht_1_90; // @[bht.scala 53:22]
  reg [1:0] pht_1_91; // @[bht.scala 53:22]
  reg [1:0] pht_1_92; // @[bht.scala 53:22]
  reg [1:0] pht_1_93; // @[bht.scala 53:22]
  reg [1:0] pht_1_94; // @[bht.scala 53:22]
  reg [1:0] pht_1_95; // @[bht.scala 53:22]
  reg [1:0] pht_1_96; // @[bht.scala 53:22]
  reg [1:0] pht_1_97; // @[bht.scala 53:22]
  reg [1:0] pht_1_98; // @[bht.scala 53:22]
  reg [1:0] pht_1_99; // @[bht.scala 53:22]
  reg [1:0] pht_1_100; // @[bht.scala 53:22]
  reg [1:0] pht_1_101; // @[bht.scala 53:22]
  reg [1:0] pht_1_102; // @[bht.scala 53:22]
  reg [1:0] pht_1_103; // @[bht.scala 53:22]
  reg [1:0] pht_1_104; // @[bht.scala 53:22]
  reg [1:0] pht_1_105; // @[bht.scala 53:22]
  reg [1:0] pht_1_106; // @[bht.scala 53:22]
  reg [1:0] pht_1_107; // @[bht.scala 53:22]
  reg [1:0] pht_1_108; // @[bht.scala 53:22]
  reg [1:0] pht_1_109; // @[bht.scala 53:22]
  reg [1:0] pht_1_110; // @[bht.scala 53:22]
  reg [1:0] pht_1_111; // @[bht.scala 53:22]
  reg [1:0] pht_1_112; // @[bht.scala 53:22]
  reg [1:0] pht_1_113; // @[bht.scala 53:22]
  reg [1:0] pht_1_114; // @[bht.scala 53:22]
  reg [1:0] pht_1_115; // @[bht.scala 53:22]
  reg [1:0] pht_1_116; // @[bht.scala 53:22]
  reg [1:0] pht_1_117; // @[bht.scala 53:22]
  reg [1:0] pht_1_118; // @[bht.scala 53:22]
  reg [1:0] pht_1_119; // @[bht.scala 53:22]
  reg [1:0] pht_1_120; // @[bht.scala 53:22]
  reg [1:0] pht_1_121; // @[bht.scala 53:22]
  reg [1:0] pht_1_122; // @[bht.scala 53:22]
  reg [1:0] pht_1_123; // @[bht.scala 53:22]
  reg [1:0] pht_1_124; // @[bht.scala 53:22]
  reg [1:0] pht_1_125; // @[bht.scala 53:22]
  reg [1:0] pht_1_126; // @[bht.scala 53:22]
  reg [1:0] pht_1_127; // @[bht.scala 53:22]
  reg [1:0] pht_1_128; // @[bht.scala 53:22]
  reg [1:0] pht_1_129; // @[bht.scala 53:22]
  reg [1:0] pht_1_130; // @[bht.scala 53:22]
  reg [1:0] pht_1_131; // @[bht.scala 53:22]
  reg [1:0] pht_1_132; // @[bht.scala 53:22]
  reg [1:0] pht_1_133; // @[bht.scala 53:22]
  reg [1:0] pht_1_134; // @[bht.scala 53:22]
  reg [1:0] pht_1_135; // @[bht.scala 53:22]
  reg [1:0] pht_1_136; // @[bht.scala 53:22]
  reg [1:0] pht_1_137; // @[bht.scala 53:22]
  reg [1:0] pht_1_138; // @[bht.scala 53:22]
  reg [1:0] pht_1_139; // @[bht.scala 53:22]
  reg [1:0] pht_1_140; // @[bht.scala 53:22]
  reg [1:0] pht_1_141; // @[bht.scala 53:22]
  reg [1:0] pht_1_142; // @[bht.scala 53:22]
  reg [1:0] pht_1_143; // @[bht.scala 53:22]
  reg [1:0] pht_1_144; // @[bht.scala 53:22]
  reg [1:0] pht_1_145; // @[bht.scala 53:22]
  reg [1:0] pht_1_146; // @[bht.scala 53:22]
  reg [1:0] pht_1_147; // @[bht.scala 53:22]
  reg [1:0] pht_1_148; // @[bht.scala 53:22]
  reg [1:0] pht_1_149; // @[bht.scala 53:22]
  reg [1:0] pht_1_150; // @[bht.scala 53:22]
  reg [1:0] pht_1_151; // @[bht.scala 53:22]
  reg [1:0] pht_1_152; // @[bht.scala 53:22]
  reg [1:0] pht_1_153; // @[bht.scala 53:22]
  reg [1:0] pht_1_154; // @[bht.scala 53:22]
  reg [1:0] pht_1_155; // @[bht.scala 53:22]
  reg [1:0] pht_1_156; // @[bht.scala 53:22]
  reg [1:0] pht_1_157; // @[bht.scala 53:22]
  reg [1:0] pht_1_158; // @[bht.scala 53:22]
  reg [1:0] pht_1_159; // @[bht.scala 53:22]
  reg [1:0] pht_1_160; // @[bht.scala 53:22]
  reg [1:0] pht_1_161; // @[bht.scala 53:22]
  reg [1:0] pht_1_162; // @[bht.scala 53:22]
  reg [1:0] pht_1_163; // @[bht.scala 53:22]
  reg [1:0] pht_1_164; // @[bht.scala 53:22]
  reg [1:0] pht_1_165; // @[bht.scala 53:22]
  reg [1:0] pht_1_166; // @[bht.scala 53:22]
  reg [1:0] pht_1_167; // @[bht.scala 53:22]
  reg [1:0] pht_1_168; // @[bht.scala 53:22]
  reg [1:0] pht_1_169; // @[bht.scala 53:22]
  reg [1:0] pht_1_170; // @[bht.scala 53:22]
  reg [1:0] pht_1_171; // @[bht.scala 53:22]
  reg [1:0] pht_1_172; // @[bht.scala 53:22]
  reg [1:0] pht_1_173; // @[bht.scala 53:22]
  reg [1:0] pht_1_174; // @[bht.scala 53:22]
  reg [1:0] pht_1_175; // @[bht.scala 53:22]
  reg [1:0] pht_1_176; // @[bht.scala 53:22]
  reg [1:0] pht_1_177; // @[bht.scala 53:22]
  reg [1:0] pht_1_178; // @[bht.scala 53:22]
  reg [1:0] pht_1_179; // @[bht.scala 53:22]
  reg [1:0] pht_1_180; // @[bht.scala 53:22]
  reg [1:0] pht_1_181; // @[bht.scala 53:22]
  reg [1:0] pht_1_182; // @[bht.scala 53:22]
  reg [1:0] pht_1_183; // @[bht.scala 53:22]
  reg [1:0] pht_1_184; // @[bht.scala 53:22]
  reg [1:0] pht_1_185; // @[bht.scala 53:22]
  reg [1:0] pht_1_186; // @[bht.scala 53:22]
  reg [1:0] pht_1_187; // @[bht.scala 53:22]
  reg [1:0] pht_1_188; // @[bht.scala 53:22]
  reg [1:0] pht_1_189; // @[bht.scala 53:22]
  reg [1:0] pht_1_190; // @[bht.scala 53:22]
  reg [1:0] pht_1_191; // @[bht.scala 53:22]
  reg [1:0] pht_1_192; // @[bht.scala 53:22]
  reg [1:0] pht_1_193; // @[bht.scala 53:22]
  reg [1:0] pht_1_194; // @[bht.scala 53:22]
  reg [1:0] pht_1_195; // @[bht.scala 53:22]
  reg [1:0] pht_1_196; // @[bht.scala 53:22]
  reg [1:0] pht_1_197; // @[bht.scala 53:22]
  reg [1:0] pht_1_198; // @[bht.scala 53:22]
  reg [1:0] pht_1_199; // @[bht.scala 53:22]
  reg [1:0] pht_1_200; // @[bht.scala 53:22]
  reg [1:0] pht_1_201; // @[bht.scala 53:22]
  reg [1:0] pht_1_202; // @[bht.scala 53:22]
  reg [1:0] pht_1_203; // @[bht.scala 53:22]
  reg [1:0] pht_1_204; // @[bht.scala 53:22]
  reg [1:0] pht_1_205; // @[bht.scala 53:22]
  reg [1:0] pht_1_206; // @[bht.scala 53:22]
  reg [1:0] pht_1_207; // @[bht.scala 53:22]
  reg [1:0] pht_1_208; // @[bht.scala 53:22]
  reg [1:0] pht_1_209; // @[bht.scala 53:22]
  reg [1:0] pht_1_210; // @[bht.scala 53:22]
  reg [1:0] pht_1_211; // @[bht.scala 53:22]
  reg [1:0] pht_1_212; // @[bht.scala 53:22]
  reg [1:0] pht_1_213; // @[bht.scala 53:22]
  reg [1:0] pht_1_214; // @[bht.scala 53:22]
  reg [1:0] pht_1_215; // @[bht.scala 53:22]
  reg [1:0] pht_1_216; // @[bht.scala 53:22]
  reg [1:0] pht_1_217; // @[bht.scala 53:22]
  reg [1:0] pht_1_218; // @[bht.scala 53:22]
  reg [1:0] pht_1_219; // @[bht.scala 53:22]
  reg [1:0] pht_1_220; // @[bht.scala 53:22]
  reg [1:0] pht_1_221; // @[bht.scala 53:22]
  reg [1:0] pht_1_222; // @[bht.scala 53:22]
  reg [1:0] pht_1_223; // @[bht.scala 53:22]
  reg [1:0] pht_1_224; // @[bht.scala 53:22]
  reg [1:0] pht_1_225; // @[bht.scala 53:22]
  reg [1:0] pht_1_226; // @[bht.scala 53:22]
  reg [1:0] pht_1_227; // @[bht.scala 53:22]
  reg [1:0] pht_1_228; // @[bht.scala 53:22]
  reg [1:0] pht_1_229; // @[bht.scala 53:22]
  reg [1:0] pht_1_230; // @[bht.scala 53:22]
  reg [1:0] pht_1_231; // @[bht.scala 53:22]
  reg [1:0] pht_1_232; // @[bht.scala 53:22]
  reg [1:0] pht_1_233; // @[bht.scala 53:22]
  reg [1:0] pht_1_234; // @[bht.scala 53:22]
  reg [1:0] pht_1_235; // @[bht.scala 53:22]
  reg [1:0] pht_1_236; // @[bht.scala 53:22]
  reg [1:0] pht_1_237; // @[bht.scala 53:22]
  reg [1:0] pht_1_238; // @[bht.scala 53:22]
  reg [1:0] pht_1_239; // @[bht.scala 53:22]
  reg [1:0] pht_1_240; // @[bht.scala 53:22]
  reg [1:0] pht_1_241; // @[bht.scala 53:22]
  reg [1:0] pht_1_242; // @[bht.scala 53:22]
  reg [1:0] pht_1_243; // @[bht.scala 53:22]
  reg [1:0] pht_1_244; // @[bht.scala 53:22]
  reg [1:0] pht_1_245; // @[bht.scala 53:22]
  reg [1:0] pht_1_246; // @[bht.scala 53:22]
  reg [1:0] pht_1_247; // @[bht.scala 53:22]
  reg [1:0] pht_1_248; // @[bht.scala 53:22]
  reg [1:0] pht_1_249; // @[bht.scala 53:22]
  reg [1:0] pht_1_250; // @[bht.scala 53:22]
  reg [1:0] pht_1_251; // @[bht.scala 53:22]
  reg [1:0] pht_1_252; // @[bht.scala 53:22]
  reg [1:0] pht_1_253; // @[bht.scala 53:22]
  reg [1:0] pht_1_254; // @[bht.scala 53:22]
  reg [1:0] pht_1_255; // @[bht.scala 53:22]
  reg [1:0] pht_2_0; // @[bht.scala 53:22]
  reg [1:0] pht_2_1; // @[bht.scala 53:22]
  reg [1:0] pht_2_2; // @[bht.scala 53:22]
  reg [1:0] pht_2_3; // @[bht.scala 53:22]
  reg [1:0] pht_2_4; // @[bht.scala 53:22]
  reg [1:0] pht_2_5; // @[bht.scala 53:22]
  reg [1:0] pht_2_6; // @[bht.scala 53:22]
  reg [1:0] pht_2_7; // @[bht.scala 53:22]
  reg [1:0] pht_2_8; // @[bht.scala 53:22]
  reg [1:0] pht_2_9; // @[bht.scala 53:22]
  reg [1:0] pht_2_10; // @[bht.scala 53:22]
  reg [1:0] pht_2_11; // @[bht.scala 53:22]
  reg [1:0] pht_2_12; // @[bht.scala 53:22]
  reg [1:0] pht_2_13; // @[bht.scala 53:22]
  reg [1:0] pht_2_14; // @[bht.scala 53:22]
  reg [1:0] pht_2_15; // @[bht.scala 53:22]
  reg [1:0] pht_2_16; // @[bht.scala 53:22]
  reg [1:0] pht_2_17; // @[bht.scala 53:22]
  reg [1:0] pht_2_18; // @[bht.scala 53:22]
  reg [1:0] pht_2_19; // @[bht.scala 53:22]
  reg [1:0] pht_2_20; // @[bht.scala 53:22]
  reg [1:0] pht_2_21; // @[bht.scala 53:22]
  reg [1:0] pht_2_22; // @[bht.scala 53:22]
  reg [1:0] pht_2_23; // @[bht.scala 53:22]
  reg [1:0] pht_2_24; // @[bht.scala 53:22]
  reg [1:0] pht_2_25; // @[bht.scala 53:22]
  reg [1:0] pht_2_26; // @[bht.scala 53:22]
  reg [1:0] pht_2_27; // @[bht.scala 53:22]
  reg [1:0] pht_2_28; // @[bht.scala 53:22]
  reg [1:0] pht_2_29; // @[bht.scala 53:22]
  reg [1:0] pht_2_30; // @[bht.scala 53:22]
  reg [1:0] pht_2_31; // @[bht.scala 53:22]
  reg [1:0] pht_2_32; // @[bht.scala 53:22]
  reg [1:0] pht_2_33; // @[bht.scala 53:22]
  reg [1:0] pht_2_34; // @[bht.scala 53:22]
  reg [1:0] pht_2_35; // @[bht.scala 53:22]
  reg [1:0] pht_2_36; // @[bht.scala 53:22]
  reg [1:0] pht_2_37; // @[bht.scala 53:22]
  reg [1:0] pht_2_38; // @[bht.scala 53:22]
  reg [1:0] pht_2_39; // @[bht.scala 53:22]
  reg [1:0] pht_2_40; // @[bht.scala 53:22]
  reg [1:0] pht_2_41; // @[bht.scala 53:22]
  reg [1:0] pht_2_42; // @[bht.scala 53:22]
  reg [1:0] pht_2_43; // @[bht.scala 53:22]
  reg [1:0] pht_2_44; // @[bht.scala 53:22]
  reg [1:0] pht_2_45; // @[bht.scala 53:22]
  reg [1:0] pht_2_46; // @[bht.scala 53:22]
  reg [1:0] pht_2_47; // @[bht.scala 53:22]
  reg [1:0] pht_2_48; // @[bht.scala 53:22]
  reg [1:0] pht_2_49; // @[bht.scala 53:22]
  reg [1:0] pht_2_50; // @[bht.scala 53:22]
  reg [1:0] pht_2_51; // @[bht.scala 53:22]
  reg [1:0] pht_2_52; // @[bht.scala 53:22]
  reg [1:0] pht_2_53; // @[bht.scala 53:22]
  reg [1:0] pht_2_54; // @[bht.scala 53:22]
  reg [1:0] pht_2_55; // @[bht.scala 53:22]
  reg [1:0] pht_2_56; // @[bht.scala 53:22]
  reg [1:0] pht_2_57; // @[bht.scala 53:22]
  reg [1:0] pht_2_58; // @[bht.scala 53:22]
  reg [1:0] pht_2_59; // @[bht.scala 53:22]
  reg [1:0] pht_2_60; // @[bht.scala 53:22]
  reg [1:0] pht_2_61; // @[bht.scala 53:22]
  reg [1:0] pht_2_62; // @[bht.scala 53:22]
  reg [1:0] pht_2_63; // @[bht.scala 53:22]
  reg [1:0] pht_2_64; // @[bht.scala 53:22]
  reg [1:0] pht_2_65; // @[bht.scala 53:22]
  reg [1:0] pht_2_66; // @[bht.scala 53:22]
  reg [1:0] pht_2_67; // @[bht.scala 53:22]
  reg [1:0] pht_2_68; // @[bht.scala 53:22]
  reg [1:0] pht_2_69; // @[bht.scala 53:22]
  reg [1:0] pht_2_70; // @[bht.scala 53:22]
  reg [1:0] pht_2_71; // @[bht.scala 53:22]
  reg [1:0] pht_2_72; // @[bht.scala 53:22]
  reg [1:0] pht_2_73; // @[bht.scala 53:22]
  reg [1:0] pht_2_74; // @[bht.scala 53:22]
  reg [1:0] pht_2_75; // @[bht.scala 53:22]
  reg [1:0] pht_2_76; // @[bht.scala 53:22]
  reg [1:0] pht_2_77; // @[bht.scala 53:22]
  reg [1:0] pht_2_78; // @[bht.scala 53:22]
  reg [1:0] pht_2_79; // @[bht.scala 53:22]
  reg [1:0] pht_2_80; // @[bht.scala 53:22]
  reg [1:0] pht_2_81; // @[bht.scala 53:22]
  reg [1:0] pht_2_82; // @[bht.scala 53:22]
  reg [1:0] pht_2_83; // @[bht.scala 53:22]
  reg [1:0] pht_2_84; // @[bht.scala 53:22]
  reg [1:0] pht_2_85; // @[bht.scala 53:22]
  reg [1:0] pht_2_86; // @[bht.scala 53:22]
  reg [1:0] pht_2_87; // @[bht.scala 53:22]
  reg [1:0] pht_2_88; // @[bht.scala 53:22]
  reg [1:0] pht_2_89; // @[bht.scala 53:22]
  reg [1:0] pht_2_90; // @[bht.scala 53:22]
  reg [1:0] pht_2_91; // @[bht.scala 53:22]
  reg [1:0] pht_2_92; // @[bht.scala 53:22]
  reg [1:0] pht_2_93; // @[bht.scala 53:22]
  reg [1:0] pht_2_94; // @[bht.scala 53:22]
  reg [1:0] pht_2_95; // @[bht.scala 53:22]
  reg [1:0] pht_2_96; // @[bht.scala 53:22]
  reg [1:0] pht_2_97; // @[bht.scala 53:22]
  reg [1:0] pht_2_98; // @[bht.scala 53:22]
  reg [1:0] pht_2_99; // @[bht.scala 53:22]
  reg [1:0] pht_2_100; // @[bht.scala 53:22]
  reg [1:0] pht_2_101; // @[bht.scala 53:22]
  reg [1:0] pht_2_102; // @[bht.scala 53:22]
  reg [1:0] pht_2_103; // @[bht.scala 53:22]
  reg [1:0] pht_2_104; // @[bht.scala 53:22]
  reg [1:0] pht_2_105; // @[bht.scala 53:22]
  reg [1:0] pht_2_106; // @[bht.scala 53:22]
  reg [1:0] pht_2_107; // @[bht.scala 53:22]
  reg [1:0] pht_2_108; // @[bht.scala 53:22]
  reg [1:0] pht_2_109; // @[bht.scala 53:22]
  reg [1:0] pht_2_110; // @[bht.scala 53:22]
  reg [1:0] pht_2_111; // @[bht.scala 53:22]
  reg [1:0] pht_2_112; // @[bht.scala 53:22]
  reg [1:0] pht_2_113; // @[bht.scala 53:22]
  reg [1:0] pht_2_114; // @[bht.scala 53:22]
  reg [1:0] pht_2_115; // @[bht.scala 53:22]
  reg [1:0] pht_2_116; // @[bht.scala 53:22]
  reg [1:0] pht_2_117; // @[bht.scala 53:22]
  reg [1:0] pht_2_118; // @[bht.scala 53:22]
  reg [1:0] pht_2_119; // @[bht.scala 53:22]
  reg [1:0] pht_2_120; // @[bht.scala 53:22]
  reg [1:0] pht_2_121; // @[bht.scala 53:22]
  reg [1:0] pht_2_122; // @[bht.scala 53:22]
  reg [1:0] pht_2_123; // @[bht.scala 53:22]
  reg [1:0] pht_2_124; // @[bht.scala 53:22]
  reg [1:0] pht_2_125; // @[bht.scala 53:22]
  reg [1:0] pht_2_126; // @[bht.scala 53:22]
  reg [1:0] pht_2_127; // @[bht.scala 53:22]
  reg [1:0] pht_2_128; // @[bht.scala 53:22]
  reg [1:0] pht_2_129; // @[bht.scala 53:22]
  reg [1:0] pht_2_130; // @[bht.scala 53:22]
  reg [1:0] pht_2_131; // @[bht.scala 53:22]
  reg [1:0] pht_2_132; // @[bht.scala 53:22]
  reg [1:0] pht_2_133; // @[bht.scala 53:22]
  reg [1:0] pht_2_134; // @[bht.scala 53:22]
  reg [1:0] pht_2_135; // @[bht.scala 53:22]
  reg [1:0] pht_2_136; // @[bht.scala 53:22]
  reg [1:0] pht_2_137; // @[bht.scala 53:22]
  reg [1:0] pht_2_138; // @[bht.scala 53:22]
  reg [1:0] pht_2_139; // @[bht.scala 53:22]
  reg [1:0] pht_2_140; // @[bht.scala 53:22]
  reg [1:0] pht_2_141; // @[bht.scala 53:22]
  reg [1:0] pht_2_142; // @[bht.scala 53:22]
  reg [1:0] pht_2_143; // @[bht.scala 53:22]
  reg [1:0] pht_2_144; // @[bht.scala 53:22]
  reg [1:0] pht_2_145; // @[bht.scala 53:22]
  reg [1:0] pht_2_146; // @[bht.scala 53:22]
  reg [1:0] pht_2_147; // @[bht.scala 53:22]
  reg [1:0] pht_2_148; // @[bht.scala 53:22]
  reg [1:0] pht_2_149; // @[bht.scala 53:22]
  reg [1:0] pht_2_150; // @[bht.scala 53:22]
  reg [1:0] pht_2_151; // @[bht.scala 53:22]
  reg [1:0] pht_2_152; // @[bht.scala 53:22]
  reg [1:0] pht_2_153; // @[bht.scala 53:22]
  reg [1:0] pht_2_154; // @[bht.scala 53:22]
  reg [1:0] pht_2_155; // @[bht.scala 53:22]
  reg [1:0] pht_2_156; // @[bht.scala 53:22]
  reg [1:0] pht_2_157; // @[bht.scala 53:22]
  reg [1:0] pht_2_158; // @[bht.scala 53:22]
  reg [1:0] pht_2_159; // @[bht.scala 53:22]
  reg [1:0] pht_2_160; // @[bht.scala 53:22]
  reg [1:0] pht_2_161; // @[bht.scala 53:22]
  reg [1:0] pht_2_162; // @[bht.scala 53:22]
  reg [1:0] pht_2_163; // @[bht.scala 53:22]
  reg [1:0] pht_2_164; // @[bht.scala 53:22]
  reg [1:0] pht_2_165; // @[bht.scala 53:22]
  reg [1:0] pht_2_166; // @[bht.scala 53:22]
  reg [1:0] pht_2_167; // @[bht.scala 53:22]
  reg [1:0] pht_2_168; // @[bht.scala 53:22]
  reg [1:0] pht_2_169; // @[bht.scala 53:22]
  reg [1:0] pht_2_170; // @[bht.scala 53:22]
  reg [1:0] pht_2_171; // @[bht.scala 53:22]
  reg [1:0] pht_2_172; // @[bht.scala 53:22]
  reg [1:0] pht_2_173; // @[bht.scala 53:22]
  reg [1:0] pht_2_174; // @[bht.scala 53:22]
  reg [1:0] pht_2_175; // @[bht.scala 53:22]
  reg [1:0] pht_2_176; // @[bht.scala 53:22]
  reg [1:0] pht_2_177; // @[bht.scala 53:22]
  reg [1:0] pht_2_178; // @[bht.scala 53:22]
  reg [1:0] pht_2_179; // @[bht.scala 53:22]
  reg [1:0] pht_2_180; // @[bht.scala 53:22]
  reg [1:0] pht_2_181; // @[bht.scala 53:22]
  reg [1:0] pht_2_182; // @[bht.scala 53:22]
  reg [1:0] pht_2_183; // @[bht.scala 53:22]
  reg [1:0] pht_2_184; // @[bht.scala 53:22]
  reg [1:0] pht_2_185; // @[bht.scala 53:22]
  reg [1:0] pht_2_186; // @[bht.scala 53:22]
  reg [1:0] pht_2_187; // @[bht.scala 53:22]
  reg [1:0] pht_2_188; // @[bht.scala 53:22]
  reg [1:0] pht_2_189; // @[bht.scala 53:22]
  reg [1:0] pht_2_190; // @[bht.scala 53:22]
  reg [1:0] pht_2_191; // @[bht.scala 53:22]
  reg [1:0] pht_2_192; // @[bht.scala 53:22]
  reg [1:0] pht_2_193; // @[bht.scala 53:22]
  reg [1:0] pht_2_194; // @[bht.scala 53:22]
  reg [1:0] pht_2_195; // @[bht.scala 53:22]
  reg [1:0] pht_2_196; // @[bht.scala 53:22]
  reg [1:0] pht_2_197; // @[bht.scala 53:22]
  reg [1:0] pht_2_198; // @[bht.scala 53:22]
  reg [1:0] pht_2_199; // @[bht.scala 53:22]
  reg [1:0] pht_2_200; // @[bht.scala 53:22]
  reg [1:0] pht_2_201; // @[bht.scala 53:22]
  reg [1:0] pht_2_202; // @[bht.scala 53:22]
  reg [1:0] pht_2_203; // @[bht.scala 53:22]
  reg [1:0] pht_2_204; // @[bht.scala 53:22]
  reg [1:0] pht_2_205; // @[bht.scala 53:22]
  reg [1:0] pht_2_206; // @[bht.scala 53:22]
  reg [1:0] pht_2_207; // @[bht.scala 53:22]
  reg [1:0] pht_2_208; // @[bht.scala 53:22]
  reg [1:0] pht_2_209; // @[bht.scala 53:22]
  reg [1:0] pht_2_210; // @[bht.scala 53:22]
  reg [1:0] pht_2_211; // @[bht.scala 53:22]
  reg [1:0] pht_2_212; // @[bht.scala 53:22]
  reg [1:0] pht_2_213; // @[bht.scala 53:22]
  reg [1:0] pht_2_214; // @[bht.scala 53:22]
  reg [1:0] pht_2_215; // @[bht.scala 53:22]
  reg [1:0] pht_2_216; // @[bht.scala 53:22]
  reg [1:0] pht_2_217; // @[bht.scala 53:22]
  reg [1:0] pht_2_218; // @[bht.scala 53:22]
  reg [1:0] pht_2_219; // @[bht.scala 53:22]
  reg [1:0] pht_2_220; // @[bht.scala 53:22]
  reg [1:0] pht_2_221; // @[bht.scala 53:22]
  reg [1:0] pht_2_222; // @[bht.scala 53:22]
  reg [1:0] pht_2_223; // @[bht.scala 53:22]
  reg [1:0] pht_2_224; // @[bht.scala 53:22]
  reg [1:0] pht_2_225; // @[bht.scala 53:22]
  reg [1:0] pht_2_226; // @[bht.scala 53:22]
  reg [1:0] pht_2_227; // @[bht.scala 53:22]
  reg [1:0] pht_2_228; // @[bht.scala 53:22]
  reg [1:0] pht_2_229; // @[bht.scala 53:22]
  reg [1:0] pht_2_230; // @[bht.scala 53:22]
  reg [1:0] pht_2_231; // @[bht.scala 53:22]
  reg [1:0] pht_2_232; // @[bht.scala 53:22]
  reg [1:0] pht_2_233; // @[bht.scala 53:22]
  reg [1:0] pht_2_234; // @[bht.scala 53:22]
  reg [1:0] pht_2_235; // @[bht.scala 53:22]
  reg [1:0] pht_2_236; // @[bht.scala 53:22]
  reg [1:0] pht_2_237; // @[bht.scala 53:22]
  reg [1:0] pht_2_238; // @[bht.scala 53:22]
  reg [1:0] pht_2_239; // @[bht.scala 53:22]
  reg [1:0] pht_2_240; // @[bht.scala 53:22]
  reg [1:0] pht_2_241; // @[bht.scala 53:22]
  reg [1:0] pht_2_242; // @[bht.scala 53:22]
  reg [1:0] pht_2_243; // @[bht.scala 53:22]
  reg [1:0] pht_2_244; // @[bht.scala 53:22]
  reg [1:0] pht_2_245; // @[bht.scala 53:22]
  reg [1:0] pht_2_246; // @[bht.scala 53:22]
  reg [1:0] pht_2_247; // @[bht.scala 53:22]
  reg [1:0] pht_2_248; // @[bht.scala 53:22]
  reg [1:0] pht_2_249; // @[bht.scala 53:22]
  reg [1:0] pht_2_250; // @[bht.scala 53:22]
  reg [1:0] pht_2_251; // @[bht.scala 53:22]
  reg [1:0] pht_2_252; // @[bht.scala 53:22]
  reg [1:0] pht_2_253; // @[bht.scala 53:22]
  reg [1:0] pht_2_254; // @[bht.scala 53:22]
  reg [1:0] pht_2_255; // @[bht.scala 53:22]
  wire [7:0] p1Addr_byte = io_pc[7:0]; // @[bht.scala 44:24]
  wire [27:0] _GEN_3329 = {{20'd0}, p1Addr_byte}; // @[bht.scala 45:22]
  wire [27:0] _p1Addr_T = 28'hce942fa ^ _GEN_3329; // @[bht.scala 45:22]
  wire [52:0] _p1Addr_T_1 = _p1Addr_T * 25'h1000193; // @[bht.scala 45:39]
  wire [7:0] p1Addr_byte_1 = io_pc[15:8]; // @[bht.scala 44:24]
  wire [52:0] _GEN_3330 = {{45'd0}, p1Addr_byte_1}; // @[bht.scala 45:22]
  wire [52:0] _p1Addr_T_2 = _p1Addr_T_1 ^ _GEN_3330; // @[bht.scala 45:22]
  wire [77:0] _p1Addr_T_3 = _p1Addr_T_2 * 25'h1000193; // @[bht.scala 45:39]
  wire [7:0] p1Addr_byte_2 = io_pc[23:16]; // @[bht.scala 44:24]
  wire [77:0] _GEN_3331 = {{70'd0}, p1Addr_byte_2}; // @[bht.scala 45:22]
  wire [77:0] _p1Addr_T_4 = _p1Addr_T_3 ^ _GEN_3331; // @[bht.scala 45:22]
  wire [102:0] _p1Addr_T_5 = _p1Addr_T_4 * 25'h1000193; // @[bht.scala 45:39]
  wire [7:0] p1Addr_byte_3 = io_pc[31:24]; // @[bht.scala 44:24]
  wire [102:0] _GEN_3332 = {{95'd0}, p1Addr_byte_3}; // @[bht.scala 45:22]
  wire [102:0] _p1Addr_T_6 = _p1Addr_T_5 ^ _GEN_3332; // @[bht.scala 45:22]
  wire [127:0] _p1Addr_T_7 = _p1Addr_T_6 * 25'h1000193; // @[bht.scala 45:39]
  wire [7:0] p1Addr = _p1Addr_T_7[7:0] ^ ghr; // @[bht.scala 50:68]
  wire [7:0] _GEN_1 = 6'h1 == _p1Addr_T_7[5:0] ? bht_1 : bht_0; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_2 = 6'h2 == _p1Addr_T_7[5:0] ? bht_2 : _GEN_1; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_3 = 6'h3 == _p1Addr_T_7[5:0] ? bht_3 : _GEN_2; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_4 = 6'h4 == _p1Addr_T_7[5:0] ? bht_4 : _GEN_3; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_5 = 6'h5 == _p1Addr_T_7[5:0] ? bht_5 : _GEN_4; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_6 = 6'h6 == _p1Addr_T_7[5:0] ? bht_6 : _GEN_5; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_7 = 6'h7 == _p1Addr_T_7[5:0] ? bht_7 : _GEN_6; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_8 = 6'h8 == _p1Addr_T_7[5:0] ? bht_8 : _GEN_7; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_9 = 6'h9 == _p1Addr_T_7[5:0] ? bht_9 : _GEN_8; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_10 = 6'ha == _p1Addr_T_7[5:0] ? bht_10 : _GEN_9; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_11 = 6'hb == _p1Addr_T_7[5:0] ? bht_11 : _GEN_10; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_12 = 6'hc == _p1Addr_T_7[5:0] ? bht_12 : _GEN_11; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_13 = 6'hd == _p1Addr_T_7[5:0] ? bht_13 : _GEN_12; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_14 = 6'he == _p1Addr_T_7[5:0] ? bht_14 : _GEN_13; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_15 = 6'hf == _p1Addr_T_7[5:0] ? bht_15 : _GEN_14; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_16 = 6'h10 == _p1Addr_T_7[5:0] ? bht_16 : _GEN_15; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_17 = 6'h11 == _p1Addr_T_7[5:0] ? bht_17 : _GEN_16; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_18 = 6'h12 == _p1Addr_T_7[5:0] ? bht_18 : _GEN_17; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_19 = 6'h13 == _p1Addr_T_7[5:0] ? bht_19 : _GEN_18; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_20 = 6'h14 == _p1Addr_T_7[5:0] ? bht_20 : _GEN_19; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_21 = 6'h15 == _p1Addr_T_7[5:0] ? bht_21 : _GEN_20; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_22 = 6'h16 == _p1Addr_T_7[5:0] ? bht_22 : _GEN_21; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_23 = 6'h17 == _p1Addr_T_7[5:0] ? bht_23 : _GEN_22; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_24 = 6'h18 == _p1Addr_T_7[5:0] ? bht_24 : _GEN_23; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_25 = 6'h19 == _p1Addr_T_7[5:0] ? bht_25 : _GEN_24; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_26 = 6'h1a == _p1Addr_T_7[5:0] ? bht_26 : _GEN_25; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_27 = 6'h1b == _p1Addr_T_7[5:0] ? bht_27 : _GEN_26; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_28 = 6'h1c == _p1Addr_T_7[5:0] ? bht_28 : _GEN_27; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_29 = 6'h1d == _p1Addr_T_7[5:0] ? bht_29 : _GEN_28; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_30 = 6'h1e == _p1Addr_T_7[5:0] ? bht_30 : _GEN_29; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_31 = 6'h1f == _p1Addr_T_7[5:0] ? bht_31 : _GEN_30; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_32 = 6'h20 == _p1Addr_T_7[5:0] ? bht_32 : _GEN_31; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_33 = 6'h21 == _p1Addr_T_7[5:0] ? bht_33 : _GEN_32; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_34 = 6'h22 == _p1Addr_T_7[5:0] ? bht_34 : _GEN_33; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_35 = 6'h23 == _p1Addr_T_7[5:0] ? bht_35 : _GEN_34; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_36 = 6'h24 == _p1Addr_T_7[5:0] ? bht_36 : _GEN_35; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_37 = 6'h25 == _p1Addr_T_7[5:0] ? bht_37 : _GEN_36; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_38 = 6'h26 == _p1Addr_T_7[5:0] ? bht_38 : _GEN_37; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_39 = 6'h27 == _p1Addr_T_7[5:0] ? bht_39 : _GEN_38; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_40 = 6'h28 == _p1Addr_T_7[5:0] ? bht_40 : _GEN_39; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_41 = 6'h29 == _p1Addr_T_7[5:0] ? bht_41 : _GEN_40; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_42 = 6'h2a == _p1Addr_T_7[5:0] ? bht_42 : _GEN_41; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_43 = 6'h2b == _p1Addr_T_7[5:0] ? bht_43 : _GEN_42; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_44 = 6'h2c == _p1Addr_T_7[5:0] ? bht_44 : _GEN_43; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_45 = 6'h2d == _p1Addr_T_7[5:0] ? bht_45 : _GEN_44; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_46 = 6'h2e == _p1Addr_T_7[5:0] ? bht_46 : _GEN_45; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_47 = 6'h2f == _p1Addr_T_7[5:0] ? bht_47 : _GEN_46; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_48 = 6'h30 == _p1Addr_T_7[5:0] ? bht_48 : _GEN_47; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_49 = 6'h31 == _p1Addr_T_7[5:0] ? bht_49 : _GEN_48; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_50 = 6'h32 == _p1Addr_T_7[5:0] ? bht_50 : _GEN_49; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_51 = 6'h33 == _p1Addr_T_7[5:0] ? bht_51 : _GEN_50; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_52 = 6'h34 == _p1Addr_T_7[5:0] ? bht_52 : _GEN_51; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_53 = 6'h35 == _p1Addr_T_7[5:0] ? bht_53 : _GEN_52; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_54 = 6'h36 == _p1Addr_T_7[5:0] ? bht_54 : _GEN_53; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_55 = 6'h37 == _p1Addr_T_7[5:0] ? bht_55 : _GEN_54; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_56 = 6'h38 == _p1Addr_T_7[5:0] ? bht_56 : _GEN_55; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_57 = 6'h39 == _p1Addr_T_7[5:0] ? bht_57 : _GEN_56; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_58 = 6'h3a == _p1Addr_T_7[5:0] ? bht_58 : _GEN_57; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_59 = 6'h3b == _p1Addr_T_7[5:0] ? bht_59 : _GEN_58; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_60 = 6'h3c == _p1Addr_T_7[5:0] ? bht_60 : _GEN_59; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_61 = 6'h3d == _p1Addr_T_7[5:0] ? bht_61 : _GEN_60; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_62 = 6'h3e == _p1Addr_T_7[5:0] ? bht_62 : _GEN_61; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_63 = 6'h3f == _p1Addr_T_7[5:0] ? bht_63 : _GEN_62; // @[bht.scala 50:{68,68}]
  wire [7:0] _pht2Data_T_9 = _p1Addr_T_7[7:0] ^ _GEN_63; // @[bht.scala 50:68]
  wire [1:0] _GEN_65 = 8'h1 == p1Addr ? pht_0_1 : pht_0_0; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_66 = 8'h2 == p1Addr ? pht_0_2 : _GEN_65; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_67 = 8'h3 == p1Addr ? pht_0_3 : _GEN_66; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_68 = 8'h4 == p1Addr ? pht_0_4 : _GEN_67; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_69 = 8'h5 == p1Addr ? pht_0_5 : _GEN_68; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_70 = 8'h6 == p1Addr ? pht_0_6 : _GEN_69; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_71 = 8'h7 == p1Addr ? pht_0_7 : _GEN_70; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_72 = 8'h8 == p1Addr ? pht_0_8 : _GEN_71; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_73 = 8'h9 == p1Addr ? pht_0_9 : _GEN_72; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_74 = 8'ha == p1Addr ? pht_0_10 : _GEN_73; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_75 = 8'hb == p1Addr ? pht_0_11 : _GEN_74; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_76 = 8'hc == p1Addr ? pht_0_12 : _GEN_75; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_77 = 8'hd == p1Addr ? pht_0_13 : _GEN_76; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_78 = 8'he == p1Addr ? pht_0_14 : _GEN_77; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_79 = 8'hf == p1Addr ? pht_0_15 : _GEN_78; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_80 = 8'h10 == p1Addr ? pht_0_16 : _GEN_79; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_81 = 8'h11 == p1Addr ? pht_0_17 : _GEN_80; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_82 = 8'h12 == p1Addr ? pht_0_18 : _GEN_81; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_83 = 8'h13 == p1Addr ? pht_0_19 : _GEN_82; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_84 = 8'h14 == p1Addr ? pht_0_20 : _GEN_83; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_85 = 8'h15 == p1Addr ? pht_0_21 : _GEN_84; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_86 = 8'h16 == p1Addr ? pht_0_22 : _GEN_85; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_87 = 8'h17 == p1Addr ? pht_0_23 : _GEN_86; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_88 = 8'h18 == p1Addr ? pht_0_24 : _GEN_87; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_89 = 8'h19 == p1Addr ? pht_0_25 : _GEN_88; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_90 = 8'h1a == p1Addr ? pht_0_26 : _GEN_89; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_91 = 8'h1b == p1Addr ? pht_0_27 : _GEN_90; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_92 = 8'h1c == p1Addr ? pht_0_28 : _GEN_91; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_93 = 8'h1d == p1Addr ? pht_0_29 : _GEN_92; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_94 = 8'h1e == p1Addr ? pht_0_30 : _GEN_93; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_95 = 8'h1f == p1Addr ? pht_0_31 : _GEN_94; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_96 = 8'h20 == p1Addr ? pht_0_32 : _GEN_95; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_97 = 8'h21 == p1Addr ? pht_0_33 : _GEN_96; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_98 = 8'h22 == p1Addr ? pht_0_34 : _GEN_97; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_99 = 8'h23 == p1Addr ? pht_0_35 : _GEN_98; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_100 = 8'h24 == p1Addr ? pht_0_36 : _GEN_99; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_101 = 8'h25 == p1Addr ? pht_0_37 : _GEN_100; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_102 = 8'h26 == p1Addr ? pht_0_38 : _GEN_101; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_103 = 8'h27 == p1Addr ? pht_0_39 : _GEN_102; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_104 = 8'h28 == p1Addr ? pht_0_40 : _GEN_103; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_105 = 8'h29 == p1Addr ? pht_0_41 : _GEN_104; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_106 = 8'h2a == p1Addr ? pht_0_42 : _GEN_105; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_107 = 8'h2b == p1Addr ? pht_0_43 : _GEN_106; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_108 = 8'h2c == p1Addr ? pht_0_44 : _GEN_107; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_109 = 8'h2d == p1Addr ? pht_0_45 : _GEN_108; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_110 = 8'h2e == p1Addr ? pht_0_46 : _GEN_109; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_111 = 8'h2f == p1Addr ? pht_0_47 : _GEN_110; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_112 = 8'h30 == p1Addr ? pht_0_48 : _GEN_111; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_113 = 8'h31 == p1Addr ? pht_0_49 : _GEN_112; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_114 = 8'h32 == p1Addr ? pht_0_50 : _GEN_113; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_115 = 8'h33 == p1Addr ? pht_0_51 : _GEN_114; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_116 = 8'h34 == p1Addr ? pht_0_52 : _GEN_115; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_117 = 8'h35 == p1Addr ? pht_0_53 : _GEN_116; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_118 = 8'h36 == p1Addr ? pht_0_54 : _GEN_117; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_119 = 8'h37 == p1Addr ? pht_0_55 : _GEN_118; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_120 = 8'h38 == p1Addr ? pht_0_56 : _GEN_119; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_121 = 8'h39 == p1Addr ? pht_0_57 : _GEN_120; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_122 = 8'h3a == p1Addr ? pht_0_58 : _GEN_121; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_123 = 8'h3b == p1Addr ? pht_0_59 : _GEN_122; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_124 = 8'h3c == p1Addr ? pht_0_60 : _GEN_123; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_125 = 8'h3d == p1Addr ? pht_0_61 : _GEN_124; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_126 = 8'h3e == p1Addr ? pht_0_62 : _GEN_125; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_127 = 8'h3f == p1Addr ? pht_0_63 : _GEN_126; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_128 = 8'h40 == p1Addr ? pht_0_64 : _GEN_127; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_129 = 8'h41 == p1Addr ? pht_0_65 : _GEN_128; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_130 = 8'h42 == p1Addr ? pht_0_66 : _GEN_129; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_131 = 8'h43 == p1Addr ? pht_0_67 : _GEN_130; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_132 = 8'h44 == p1Addr ? pht_0_68 : _GEN_131; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_133 = 8'h45 == p1Addr ? pht_0_69 : _GEN_132; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_134 = 8'h46 == p1Addr ? pht_0_70 : _GEN_133; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_135 = 8'h47 == p1Addr ? pht_0_71 : _GEN_134; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_136 = 8'h48 == p1Addr ? pht_0_72 : _GEN_135; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_137 = 8'h49 == p1Addr ? pht_0_73 : _GEN_136; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_138 = 8'h4a == p1Addr ? pht_0_74 : _GEN_137; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_139 = 8'h4b == p1Addr ? pht_0_75 : _GEN_138; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_140 = 8'h4c == p1Addr ? pht_0_76 : _GEN_139; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_141 = 8'h4d == p1Addr ? pht_0_77 : _GEN_140; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_142 = 8'h4e == p1Addr ? pht_0_78 : _GEN_141; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_143 = 8'h4f == p1Addr ? pht_0_79 : _GEN_142; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_144 = 8'h50 == p1Addr ? pht_0_80 : _GEN_143; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_145 = 8'h51 == p1Addr ? pht_0_81 : _GEN_144; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_146 = 8'h52 == p1Addr ? pht_0_82 : _GEN_145; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_147 = 8'h53 == p1Addr ? pht_0_83 : _GEN_146; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_148 = 8'h54 == p1Addr ? pht_0_84 : _GEN_147; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_149 = 8'h55 == p1Addr ? pht_0_85 : _GEN_148; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_150 = 8'h56 == p1Addr ? pht_0_86 : _GEN_149; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_151 = 8'h57 == p1Addr ? pht_0_87 : _GEN_150; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_152 = 8'h58 == p1Addr ? pht_0_88 : _GEN_151; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_153 = 8'h59 == p1Addr ? pht_0_89 : _GEN_152; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_154 = 8'h5a == p1Addr ? pht_0_90 : _GEN_153; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_155 = 8'h5b == p1Addr ? pht_0_91 : _GEN_154; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_156 = 8'h5c == p1Addr ? pht_0_92 : _GEN_155; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_157 = 8'h5d == p1Addr ? pht_0_93 : _GEN_156; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_158 = 8'h5e == p1Addr ? pht_0_94 : _GEN_157; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_159 = 8'h5f == p1Addr ? pht_0_95 : _GEN_158; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_160 = 8'h60 == p1Addr ? pht_0_96 : _GEN_159; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_161 = 8'h61 == p1Addr ? pht_0_97 : _GEN_160; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_162 = 8'h62 == p1Addr ? pht_0_98 : _GEN_161; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_163 = 8'h63 == p1Addr ? pht_0_99 : _GEN_162; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_164 = 8'h64 == p1Addr ? pht_0_100 : _GEN_163; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_165 = 8'h65 == p1Addr ? pht_0_101 : _GEN_164; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_166 = 8'h66 == p1Addr ? pht_0_102 : _GEN_165; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_167 = 8'h67 == p1Addr ? pht_0_103 : _GEN_166; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_168 = 8'h68 == p1Addr ? pht_0_104 : _GEN_167; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_169 = 8'h69 == p1Addr ? pht_0_105 : _GEN_168; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_170 = 8'h6a == p1Addr ? pht_0_106 : _GEN_169; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_171 = 8'h6b == p1Addr ? pht_0_107 : _GEN_170; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_172 = 8'h6c == p1Addr ? pht_0_108 : _GEN_171; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_173 = 8'h6d == p1Addr ? pht_0_109 : _GEN_172; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_174 = 8'h6e == p1Addr ? pht_0_110 : _GEN_173; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_175 = 8'h6f == p1Addr ? pht_0_111 : _GEN_174; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_176 = 8'h70 == p1Addr ? pht_0_112 : _GEN_175; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_177 = 8'h71 == p1Addr ? pht_0_113 : _GEN_176; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_178 = 8'h72 == p1Addr ? pht_0_114 : _GEN_177; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_179 = 8'h73 == p1Addr ? pht_0_115 : _GEN_178; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_180 = 8'h74 == p1Addr ? pht_0_116 : _GEN_179; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_181 = 8'h75 == p1Addr ? pht_0_117 : _GEN_180; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_182 = 8'h76 == p1Addr ? pht_0_118 : _GEN_181; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_183 = 8'h77 == p1Addr ? pht_0_119 : _GEN_182; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_184 = 8'h78 == p1Addr ? pht_0_120 : _GEN_183; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_185 = 8'h79 == p1Addr ? pht_0_121 : _GEN_184; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_186 = 8'h7a == p1Addr ? pht_0_122 : _GEN_185; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_187 = 8'h7b == p1Addr ? pht_0_123 : _GEN_186; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_188 = 8'h7c == p1Addr ? pht_0_124 : _GEN_187; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_189 = 8'h7d == p1Addr ? pht_0_125 : _GEN_188; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_190 = 8'h7e == p1Addr ? pht_0_126 : _GEN_189; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_191 = 8'h7f == p1Addr ? pht_0_127 : _GEN_190; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_192 = 8'h80 == p1Addr ? pht_0_128 : _GEN_191; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_193 = 8'h81 == p1Addr ? pht_0_129 : _GEN_192; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_194 = 8'h82 == p1Addr ? pht_0_130 : _GEN_193; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_195 = 8'h83 == p1Addr ? pht_0_131 : _GEN_194; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_196 = 8'h84 == p1Addr ? pht_0_132 : _GEN_195; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_197 = 8'h85 == p1Addr ? pht_0_133 : _GEN_196; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_198 = 8'h86 == p1Addr ? pht_0_134 : _GEN_197; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_199 = 8'h87 == p1Addr ? pht_0_135 : _GEN_198; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_200 = 8'h88 == p1Addr ? pht_0_136 : _GEN_199; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_201 = 8'h89 == p1Addr ? pht_0_137 : _GEN_200; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_202 = 8'h8a == p1Addr ? pht_0_138 : _GEN_201; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_203 = 8'h8b == p1Addr ? pht_0_139 : _GEN_202; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_204 = 8'h8c == p1Addr ? pht_0_140 : _GEN_203; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_205 = 8'h8d == p1Addr ? pht_0_141 : _GEN_204; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_206 = 8'h8e == p1Addr ? pht_0_142 : _GEN_205; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_207 = 8'h8f == p1Addr ? pht_0_143 : _GEN_206; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_208 = 8'h90 == p1Addr ? pht_0_144 : _GEN_207; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_209 = 8'h91 == p1Addr ? pht_0_145 : _GEN_208; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_210 = 8'h92 == p1Addr ? pht_0_146 : _GEN_209; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_211 = 8'h93 == p1Addr ? pht_0_147 : _GEN_210; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_212 = 8'h94 == p1Addr ? pht_0_148 : _GEN_211; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_213 = 8'h95 == p1Addr ? pht_0_149 : _GEN_212; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_214 = 8'h96 == p1Addr ? pht_0_150 : _GEN_213; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_215 = 8'h97 == p1Addr ? pht_0_151 : _GEN_214; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_216 = 8'h98 == p1Addr ? pht_0_152 : _GEN_215; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_217 = 8'h99 == p1Addr ? pht_0_153 : _GEN_216; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_218 = 8'h9a == p1Addr ? pht_0_154 : _GEN_217; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_219 = 8'h9b == p1Addr ? pht_0_155 : _GEN_218; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_220 = 8'h9c == p1Addr ? pht_0_156 : _GEN_219; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_221 = 8'h9d == p1Addr ? pht_0_157 : _GEN_220; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_222 = 8'h9e == p1Addr ? pht_0_158 : _GEN_221; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_223 = 8'h9f == p1Addr ? pht_0_159 : _GEN_222; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_224 = 8'ha0 == p1Addr ? pht_0_160 : _GEN_223; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_225 = 8'ha1 == p1Addr ? pht_0_161 : _GEN_224; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_226 = 8'ha2 == p1Addr ? pht_0_162 : _GEN_225; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_227 = 8'ha3 == p1Addr ? pht_0_163 : _GEN_226; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_228 = 8'ha4 == p1Addr ? pht_0_164 : _GEN_227; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_229 = 8'ha5 == p1Addr ? pht_0_165 : _GEN_228; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_230 = 8'ha6 == p1Addr ? pht_0_166 : _GEN_229; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_231 = 8'ha7 == p1Addr ? pht_0_167 : _GEN_230; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_232 = 8'ha8 == p1Addr ? pht_0_168 : _GEN_231; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_233 = 8'ha9 == p1Addr ? pht_0_169 : _GEN_232; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_234 = 8'haa == p1Addr ? pht_0_170 : _GEN_233; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_235 = 8'hab == p1Addr ? pht_0_171 : _GEN_234; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_236 = 8'hac == p1Addr ? pht_0_172 : _GEN_235; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_237 = 8'had == p1Addr ? pht_0_173 : _GEN_236; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_238 = 8'hae == p1Addr ? pht_0_174 : _GEN_237; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_239 = 8'haf == p1Addr ? pht_0_175 : _GEN_238; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_240 = 8'hb0 == p1Addr ? pht_0_176 : _GEN_239; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_241 = 8'hb1 == p1Addr ? pht_0_177 : _GEN_240; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_242 = 8'hb2 == p1Addr ? pht_0_178 : _GEN_241; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_243 = 8'hb3 == p1Addr ? pht_0_179 : _GEN_242; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_244 = 8'hb4 == p1Addr ? pht_0_180 : _GEN_243; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_245 = 8'hb5 == p1Addr ? pht_0_181 : _GEN_244; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_246 = 8'hb6 == p1Addr ? pht_0_182 : _GEN_245; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_247 = 8'hb7 == p1Addr ? pht_0_183 : _GEN_246; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_248 = 8'hb8 == p1Addr ? pht_0_184 : _GEN_247; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_249 = 8'hb9 == p1Addr ? pht_0_185 : _GEN_248; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_250 = 8'hba == p1Addr ? pht_0_186 : _GEN_249; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_251 = 8'hbb == p1Addr ? pht_0_187 : _GEN_250; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_252 = 8'hbc == p1Addr ? pht_0_188 : _GEN_251; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_253 = 8'hbd == p1Addr ? pht_0_189 : _GEN_252; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_254 = 8'hbe == p1Addr ? pht_0_190 : _GEN_253; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_255 = 8'hbf == p1Addr ? pht_0_191 : _GEN_254; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_256 = 8'hc0 == p1Addr ? pht_0_192 : _GEN_255; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_257 = 8'hc1 == p1Addr ? pht_0_193 : _GEN_256; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_258 = 8'hc2 == p1Addr ? pht_0_194 : _GEN_257; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_259 = 8'hc3 == p1Addr ? pht_0_195 : _GEN_258; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_260 = 8'hc4 == p1Addr ? pht_0_196 : _GEN_259; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_261 = 8'hc5 == p1Addr ? pht_0_197 : _GEN_260; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_262 = 8'hc6 == p1Addr ? pht_0_198 : _GEN_261; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_263 = 8'hc7 == p1Addr ? pht_0_199 : _GEN_262; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_264 = 8'hc8 == p1Addr ? pht_0_200 : _GEN_263; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_265 = 8'hc9 == p1Addr ? pht_0_201 : _GEN_264; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_266 = 8'hca == p1Addr ? pht_0_202 : _GEN_265; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_267 = 8'hcb == p1Addr ? pht_0_203 : _GEN_266; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_268 = 8'hcc == p1Addr ? pht_0_204 : _GEN_267; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_269 = 8'hcd == p1Addr ? pht_0_205 : _GEN_268; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_270 = 8'hce == p1Addr ? pht_0_206 : _GEN_269; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_271 = 8'hcf == p1Addr ? pht_0_207 : _GEN_270; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_272 = 8'hd0 == p1Addr ? pht_0_208 : _GEN_271; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_273 = 8'hd1 == p1Addr ? pht_0_209 : _GEN_272; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_274 = 8'hd2 == p1Addr ? pht_0_210 : _GEN_273; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_275 = 8'hd3 == p1Addr ? pht_0_211 : _GEN_274; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_276 = 8'hd4 == p1Addr ? pht_0_212 : _GEN_275; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_277 = 8'hd5 == p1Addr ? pht_0_213 : _GEN_276; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_278 = 8'hd6 == p1Addr ? pht_0_214 : _GEN_277; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_279 = 8'hd7 == p1Addr ? pht_0_215 : _GEN_278; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_280 = 8'hd8 == p1Addr ? pht_0_216 : _GEN_279; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_281 = 8'hd9 == p1Addr ? pht_0_217 : _GEN_280; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_282 = 8'hda == p1Addr ? pht_0_218 : _GEN_281; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_283 = 8'hdb == p1Addr ? pht_0_219 : _GEN_282; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_284 = 8'hdc == p1Addr ? pht_0_220 : _GEN_283; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_285 = 8'hdd == p1Addr ? pht_0_221 : _GEN_284; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_286 = 8'hde == p1Addr ? pht_0_222 : _GEN_285; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_287 = 8'hdf == p1Addr ? pht_0_223 : _GEN_286; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_288 = 8'he0 == p1Addr ? pht_0_224 : _GEN_287; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_289 = 8'he1 == p1Addr ? pht_0_225 : _GEN_288; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_290 = 8'he2 == p1Addr ? pht_0_226 : _GEN_289; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_291 = 8'he3 == p1Addr ? pht_0_227 : _GEN_290; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_292 = 8'he4 == p1Addr ? pht_0_228 : _GEN_291; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_293 = 8'he5 == p1Addr ? pht_0_229 : _GEN_292; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_294 = 8'he6 == p1Addr ? pht_0_230 : _GEN_293; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_295 = 8'he7 == p1Addr ? pht_0_231 : _GEN_294; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_296 = 8'he8 == p1Addr ? pht_0_232 : _GEN_295; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_297 = 8'he9 == p1Addr ? pht_0_233 : _GEN_296; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_298 = 8'hea == p1Addr ? pht_0_234 : _GEN_297; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_299 = 8'heb == p1Addr ? pht_0_235 : _GEN_298; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_300 = 8'hec == p1Addr ? pht_0_236 : _GEN_299; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_301 = 8'hed == p1Addr ? pht_0_237 : _GEN_300; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_302 = 8'hee == p1Addr ? pht_0_238 : _GEN_301; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_303 = 8'hef == p1Addr ? pht_0_239 : _GEN_302; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_304 = 8'hf0 == p1Addr ? pht_0_240 : _GEN_303; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_305 = 8'hf1 == p1Addr ? pht_0_241 : _GEN_304; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_306 = 8'hf2 == p1Addr ? pht_0_242 : _GEN_305; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_307 = 8'hf3 == p1Addr ? pht_0_243 : _GEN_306; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_308 = 8'hf4 == p1Addr ? pht_0_244 : _GEN_307; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_309 = 8'hf5 == p1Addr ? pht_0_245 : _GEN_308; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_310 = 8'hf6 == p1Addr ? pht_0_246 : _GEN_309; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_311 = 8'hf7 == p1Addr ? pht_0_247 : _GEN_310; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_312 = 8'hf8 == p1Addr ? pht_0_248 : _GEN_311; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_313 = 8'hf9 == p1Addr ? pht_0_249 : _GEN_312; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_314 = 8'hfa == p1Addr ? pht_0_250 : _GEN_313; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_315 = 8'hfb == p1Addr ? pht_0_251 : _GEN_314; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_316 = 8'hfc == p1Addr ? pht_0_252 : _GEN_315; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_317 = 8'hfd == p1Addr ? pht_0_253 : _GEN_316; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_318 = 8'hfe == p1Addr ? pht_0_254 : _GEN_317; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_319 = 8'hff == p1Addr ? pht_0_255 : _GEN_318; // @[bht.scala 60:{32,32}]
  wire [1:0] _GEN_321 = 8'h1 == _pht2Data_T_9 ? pht_2_1 : pht_2_0; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_322 = 8'h2 == _pht2Data_T_9 ? pht_2_2 : _GEN_321; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_323 = 8'h3 == _pht2Data_T_9 ? pht_2_3 : _GEN_322; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_324 = 8'h4 == _pht2Data_T_9 ? pht_2_4 : _GEN_323; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_325 = 8'h5 == _pht2Data_T_9 ? pht_2_5 : _GEN_324; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_326 = 8'h6 == _pht2Data_T_9 ? pht_2_6 : _GEN_325; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_327 = 8'h7 == _pht2Data_T_9 ? pht_2_7 : _GEN_326; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_328 = 8'h8 == _pht2Data_T_9 ? pht_2_8 : _GEN_327; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_329 = 8'h9 == _pht2Data_T_9 ? pht_2_9 : _GEN_328; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_330 = 8'ha == _pht2Data_T_9 ? pht_2_10 : _GEN_329; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_331 = 8'hb == _pht2Data_T_9 ? pht_2_11 : _GEN_330; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_332 = 8'hc == _pht2Data_T_9 ? pht_2_12 : _GEN_331; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_333 = 8'hd == _pht2Data_T_9 ? pht_2_13 : _GEN_332; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_334 = 8'he == _pht2Data_T_9 ? pht_2_14 : _GEN_333; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_335 = 8'hf == _pht2Data_T_9 ? pht_2_15 : _GEN_334; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_336 = 8'h10 == _pht2Data_T_9 ? pht_2_16 : _GEN_335; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_337 = 8'h11 == _pht2Data_T_9 ? pht_2_17 : _GEN_336; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_338 = 8'h12 == _pht2Data_T_9 ? pht_2_18 : _GEN_337; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_339 = 8'h13 == _pht2Data_T_9 ? pht_2_19 : _GEN_338; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_340 = 8'h14 == _pht2Data_T_9 ? pht_2_20 : _GEN_339; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_341 = 8'h15 == _pht2Data_T_9 ? pht_2_21 : _GEN_340; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_342 = 8'h16 == _pht2Data_T_9 ? pht_2_22 : _GEN_341; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_343 = 8'h17 == _pht2Data_T_9 ? pht_2_23 : _GEN_342; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_344 = 8'h18 == _pht2Data_T_9 ? pht_2_24 : _GEN_343; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_345 = 8'h19 == _pht2Data_T_9 ? pht_2_25 : _GEN_344; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_346 = 8'h1a == _pht2Data_T_9 ? pht_2_26 : _GEN_345; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_347 = 8'h1b == _pht2Data_T_9 ? pht_2_27 : _GEN_346; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_348 = 8'h1c == _pht2Data_T_9 ? pht_2_28 : _GEN_347; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_349 = 8'h1d == _pht2Data_T_9 ? pht_2_29 : _GEN_348; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_350 = 8'h1e == _pht2Data_T_9 ? pht_2_30 : _GEN_349; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_351 = 8'h1f == _pht2Data_T_9 ? pht_2_31 : _GEN_350; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_352 = 8'h20 == _pht2Data_T_9 ? pht_2_32 : _GEN_351; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_353 = 8'h21 == _pht2Data_T_9 ? pht_2_33 : _GEN_352; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_354 = 8'h22 == _pht2Data_T_9 ? pht_2_34 : _GEN_353; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_355 = 8'h23 == _pht2Data_T_9 ? pht_2_35 : _GEN_354; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_356 = 8'h24 == _pht2Data_T_9 ? pht_2_36 : _GEN_355; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_357 = 8'h25 == _pht2Data_T_9 ? pht_2_37 : _GEN_356; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_358 = 8'h26 == _pht2Data_T_9 ? pht_2_38 : _GEN_357; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_359 = 8'h27 == _pht2Data_T_9 ? pht_2_39 : _GEN_358; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_360 = 8'h28 == _pht2Data_T_9 ? pht_2_40 : _GEN_359; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_361 = 8'h29 == _pht2Data_T_9 ? pht_2_41 : _GEN_360; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_362 = 8'h2a == _pht2Data_T_9 ? pht_2_42 : _GEN_361; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_363 = 8'h2b == _pht2Data_T_9 ? pht_2_43 : _GEN_362; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_364 = 8'h2c == _pht2Data_T_9 ? pht_2_44 : _GEN_363; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_365 = 8'h2d == _pht2Data_T_9 ? pht_2_45 : _GEN_364; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_366 = 8'h2e == _pht2Data_T_9 ? pht_2_46 : _GEN_365; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_367 = 8'h2f == _pht2Data_T_9 ? pht_2_47 : _GEN_366; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_368 = 8'h30 == _pht2Data_T_9 ? pht_2_48 : _GEN_367; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_369 = 8'h31 == _pht2Data_T_9 ? pht_2_49 : _GEN_368; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_370 = 8'h32 == _pht2Data_T_9 ? pht_2_50 : _GEN_369; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_371 = 8'h33 == _pht2Data_T_9 ? pht_2_51 : _GEN_370; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_372 = 8'h34 == _pht2Data_T_9 ? pht_2_52 : _GEN_371; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_373 = 8'h35 == _pht2Data_T_9 ? pht_2_53 : _GEN_372; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_374 = 8'h36 == _pht2Data_T_9 ? pht_2_54 : _GEN_373; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_375 = 8'h37 == _pht2Data_T_9 ? pht_2_55 : _GEN_374; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_376 = 8'h38 == _pht2Data_T_9 ? pht_2_56 : _GEN_375; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_377 = 8'h39 == _pht2Data_T_9 ? pht_2_57 : _GEN_376; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_378 = 8'h3a == _pht2Data_T_9 ? pht_2_58 : _GEN_377; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_379 = 8'h3b == _pht2Data_T_9 ? pht_2_59 : _GEN_378; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_380 = 8'h3c == _pht2Data_T_9 ? pht_2_60 : _GEN_379; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_381 = 8'h3d == _pht2Data_T_9 ? pht_2_61 : _GEN_380; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_382 = 8'h3e == _pht2Data_T_9 ? pht_2_62 : _GEN_381; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_383 = 8'h3f == _pht2Data_T_9 ? pht_2_63 : _GEN_382; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_384 = 8'h40 == _pht2Data_T_9 ? pht_2_64 : _GEN_383; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_385 = 8'h41 == _pht2Data_T_9 ? pht_2_65 : _GEN_384; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_386 = 8'h42 == _pht2Data_T_9 ? pht_2_66 : _GEN_385; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_387 = 8'h43 == _pht2Data_T_9 ? pht_2_67 : _GEN_386; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_388 = 8'h44 == _pht2Data_T_9 ? pht_2_68 : _GEN_387; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_389 = 8'h45 == _pht2Data_T_9 ? pht_2_69 : _GEN_388; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_390 = 8'h46 == _pht2Data_T_9 ? pht_2_70 : _GEN_389; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_391 = 8'h47 == _pht2Data_T_9 ? pht_2_71 : _GEN_390; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_392 = 8'h48 == _pht2Data_T_9 ? pht_2_72 : _GEN_391; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_393 = 8'h49 == _pht2Data_T_9 ? pht_2_73 : _GEN_392; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_394 = 8'h4a == _pht2Data_T_9 ? pht_2_74 : _GEN_393; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_395 = 8'h4b == _pht2Data_T_9 ? pht_2_75 : _GEN_394; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_396 = 8'h4c == _pht2Data_T_9 ? pht_2_76 : _GEN_395; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_397 = 8'h4d == _pht2Data_T_9 ? pht_2_77 : _GEN_396; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_398 = 8'h4e == _pht2Data_T_9 ? pht_2_78 : _GEN_397; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_399 = 8'h4f == _pht2Data_T_9 ? pht_2_79 : _GEN_398; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_400 = 8'h50 == _pht2Data_T_9 ? pht_2_80 : _GEN_399; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_401 = 8'h51 == _pht2Data_T_9 ? pht_2_81 : _GEN_400; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_402 = 8'h52 == _pht2Data_T_9 ? pht_2_82 : _GEN_401; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_403 = 8'h53 == _pht2Data_T_9 ? pht_2_83 : _GEN_402; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_404 = 8'h54 == _pht2Data_T_9 ? pht_2_84 : _GEN_403; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_405 = 8'h55 == _pht2Data_T_9 ? pht_2_85 : _GEN_404; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_406 = 8'h56 == _pht2Data_T_9 ? pht_2_86 : _GEN_405; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_407 = 8'h57 == _pht2Data_T_9 ? pht_2_87 : _GEN_406; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_408 = 8'h58 == _pht2Data_T_9 ? pht_2_88 : _GEN_407; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_409 = 8'h59 == _pht2Data_T_9 ? pht_2_89 : _GEN_408; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_410 = 8'h5a == _pht2Data_T_9 ? pht_2_90 : _GEN_409; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_411 = 8'h5b == _pht2Data_T_9 ? pht_2_91 : _GEN_410; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_412 = 8'h5c == _pht2Data_T_9 ? pht_2_92 : _GEN_411; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_413 = 8'h5d == _pht2Data_T_9 ? pht_2_93 : _GEN_412; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_414 = 8'h5e == _pht2Data_T_9 ? pht_2_94 : _GEN_413; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_415 = 8'h5f == _pht2Data_T_9 ? pht_2_95 : _GEN_414; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_416 = 8'h60 == _pht2Data_T_9 ? pht_2_96 : _GEN_415; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_417 = 8'h61 == _pht2Data_T_9 ? pht_2_97 : _GEN_416; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_418 = 8'h62 == _pht2Data_T_9 ? pht_2_98 : _GEN_417; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_419 = 8'h63 == _pht2Data_T_9 ? pht_2_99 : _GEN_418; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_420 = 8'h64 == _pht2Data_T_9 ? pht_2_100 : _GEN_419; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_421 = 8'h65 == _pht2Data_T_9 ? pht_2_101 : _GEN_420; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_422 = 8'h66 == _pht2Data_T_9 ? pht_2_102 : _GEN_421; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_423 = 8'h67 == _pht2Data_T_9 ? pht_2_103 : _GEN_422; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_424 = 8'h68 == _pht2Data_T_9 ? pht_2_104 : _GEN_423; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_425 = 8'h69 == _pht2Data_T_9 ? pht_2_105 : _GEN_424; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_426 = 8'h6a == _pht2Data_T_9 ? pht_2_106 : _GEN_425; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_427 = 8'h6b == _pht2Data_T_9 ? pht_2_107 : _GEN_426; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_428 = 8'h6c == _pht2Data_T_9 ? pht_2_108 : _GEN_427; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_429 = 8'h6d == _pht2Data_T_9 ? pht_2_109 : _GEN_428; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_430 = 8'h6e == _pht2Data_T_9 ? pht_2_110 : _GEN_429; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_431 = 8'h6f == _pht2Data_T_9 ? pht_2_111 : _GEN_430; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_432 = 8'h70 == _pht2Data_T_9 ? pht_2_112 : _GEN_431; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_433 = 8'h71 == _pht2Data_T_9 ? pht_2_113 : _GEN_432; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_434 = 8'h72 == _pht2Data_T_9 ? pht_2_114 : _GEN_433; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_435 = 8'h73 == _pht2Data_T_9 ? pht_2_115 : _GEN_434; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_436 = 8'h74 == _pht2Data_T_9 ? pht_2_116 : _GEN_435; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_437 = 8'h75 == _pht2Data_T_9 ? pht_2_117 : _GEN_436; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_438 = 8'h76 == _pht2Data_T_9 ? pht_2_118 : _GEN_437; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_439 = 8'h77 == _pht2Data_T_9 ? pht_2_119 : _GEN_438; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_440 = 8'h78 == _pht2Data_T_9 ? pht_2_120 : _GEN_439; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_441 = 8'h79 == _pht2Data_T_9 ? pht_2_121 : _GEN_440; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_442 = 8'h7a == _pht2Data_T_9 ? pht_2_122 : _GEN_441; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_443 = 8'h7b == _pht2Data_T_9 ? pht_2_123 : _GEN_442; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_444 = 8'h7c == _pht2Data_T_9 ? pht_2_124 : _GEN_443; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_445 = 8'h7d == _pht2Data_T_9 ? pht_2_125 : _GEN_444; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_446 = 8'h7e == _pht2Data_T_9 ? pht_2_126 : _GEN_445; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_447 = 8'h7f == _pht2Data_T_9 ? pht_2_127 : _GEN_446; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_448 = 8'h80 == _pht2Data_T_9 ? pht_2_128 : _GEN_447; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_449 = 8'h81 == _pht2Data_T_9 ? pht_2_129 : _GEN_448; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_450 = 8'h82 == _pht2Data_T_9 ? pht_2_130 : _GEN_449; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_451 = 8'h83 == _pht2Data_T_9 ? pht_2_131 : _GEN_450; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_452 = 8'h84 == _pht2Data_T_9 ? pht_2_132 : _GEN_451; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_453 = 8'h85 == _pht2Data_T_9 ? pht_2_133 : _GEN_452; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_454 = 8'h86 == _pht2Data_T_9 ? pht_2_134 : _GEN_453; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_455 = 8'h87 == _pht2Data_T_9 ? pht_2_135 : _GEN_454; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_456 = 8'h88 == _pht2Data_T_9 ? pht_2_136 : _GEN_455; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_457 = 8'h89 == _pht2Data_T_9 ? pht_2_137 : _GEN_456; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_458 = 8'h8a == _pht2Data_T_9 ? pht_2_138 : _GEN_457; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_459 = 8'h8b == _pht2Data_T_9 ? pht_2_139 : _GEN_458; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_460 = 8'h8c == _pht2Data_T_9 ? pht_2_140 : _GEN_459; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_461 = 8'h8d == _pht2Data_T_9 ? pht_2_141 : _GEN_460; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_462 = 8'h8e == _pht2Data_T_9 ? pht_2_142 : _GEN_461; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_463 = 8'h8f == _pht2Data_T_9 ? pht_2_143 : _GEN_462; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_464 = 8'h90 == _pht2Data_T_9 ? pht_2_144 : _GEN_463; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_465 = 8'h91 == _pht2Data_T_9 ? pht_2_145 : _GEN_464; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_466 = 8'h92 == _pht2Data_T_9 ? pht_2_146 : _GEN_465; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_467 = 8'h93 == _pht2Data_T_9 ? pht_2_147 : _GEN_466; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_468 = 8'h94 == _pht2Data_T_9 ? pht_2_148 : _GEN_467; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_469 = 8'h95 == _pht2Data_T_9 ? pht_2_149 : _GEN_468; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_470 = 8'h96 == _pht2Data_T_9 ? pht_2_150 : _GEN_469; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_471 = 8'h97 == _pht2Data_T_9 ? pht_2_151 : _GEN_470; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_472 = 8'h98 == _pht2Data_T_9 ? pht_2_152 : _GEN_471; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_473 = 8'h99 == _pht2Data_T_9 ? pht_2_153 : _GEN_472; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_474 = 8'h9a == _pht2Data_T_9 ? pht_2_154 : _GEN_473; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_475 = 8'h9b == _pht2Data_T_9 ? pht_2_155 : _GEN_474; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_476 = 8'h9c == _pht2Data_T_9 ? pht_2_156 : _GEN_475; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_477 = 8'h9d == _pht2Data_T_9 ? pht_2_157 : _GEN_476; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_478 = 8'h9e == _pht2Data_T_9 ? pht_2_158 : _GEN_477; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_479 = 8'h9f == _pht2Data_T_9 ? pht_2_159 : _GEN_478; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_480 = 8'ha0 == _pht2Data_T_9 ? pht_2_160 : _GEN_479; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_481 = 8'ha1 == _pht2Data_T_9 ? pht_2_161 : _GEN_480; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_482 = 8'ha2 == _pht2Data_T_9 ? pht_2_162 : _GEN_481; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_483 = 8'ha3 == _pht2Data_T_9 ? pht_2_163 : _GEN_482; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_484 = 8'ha4 == _pht2Data_T_9 ? pht_2_164 : _GEN_483; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_485 = 8'ha5 == _pht2Data_T_9 ? pht_2_165 : _GEN_484; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_486 = 8'ha6 == _pht2Data_T_9 ? pht_2_166 : _GEN_485; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_487 = 8'ha7 == _pht2Data_T_9 ? pht_2_167 : _GEN_486; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_488 = 8'ha8 == _pht2Data_T_9 ? pht_2_168 : _GEN_487; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_489 = 8'ha9 == _pht2Data_T_9 ? pht_2_169 : _GEN_488; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_490 = 8'haa == _pht2Data_T_9 ? pht_2_170 : _GEN_489; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_491 = 8'hab == _pht2Data_T_9 ? pht_2_171 : _GEN_490; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_492 = 8'hac == _pht2Data_T_9 ? pht_2_172 : _GEN_491; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_493 = 8'had == _pht2Data_T_9 ? pht_2_173 : _GEN_492; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_494 = 8'hae == _pht2Data_T_9 ? pht_2_174 : _GEN_493; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_495 = 8'haf == _pht2Data_T_9 ? pht_2_175 : _GEN_494; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_496 = 8'hb0 == _pht2Data_T_9 ? pht_2_176 : _GEN_495; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_497 = 8'hb1 == _pht2Data_T_9 ? pht_2_177 : _GEN_496; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_498 = 8'hb2 == _pht2Data_T_9 ? pht_2_178 : _GEN_497; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_499 = 8'hb3 == _pht2Data_T_9 ? pht_2_179 : _GEN_498; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_500 = 8'hb4 == _pht2Data_T_9 ? pht_2_180 : _GEN_499; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_501 = 8'hb5 == _pht2Data_T_9 ? pht_2_181 : _GEN_500; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_502 = 8'hb6 == _pht2Data_T_9 ? pht_2_182 : _GEN_501; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_503 = 8'hb7 == _pht2Data_T_9 ? pht_2_183 : _GEN_502; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_504 = 8'hb8 == _pht2Data_T_9 ? pht_2_184 : _GEN_503; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_505 = 8'hb9 == _pht2Data_T_9 ? pht_2_185 : _GEN_504; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_506 = 8'hba == _pht2Data_T_9 ? pht_2_186 : _GEN_505; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_507 = 8'hbb == _pht2Data_T_9 ? pht_2_187 : _GEN_506; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_508 = 8'hbc == _pht2Data_T_9 ? pht_2_188 : _GEN_507; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_509 = 8'hbd == _pht2Data_T_9 ? pht_2_189 : _GEN_508; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_510 = 8'hbe == _pht2Data_T_9 ? pht_2_190 : _GEN_509; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_511 = 8'hbf == _pht2Data_T_9 ? pht_2_191 : _GEN_510; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_512 = 8'hc0 == _pht2Data_T_9 ? pht_2_192 : _GEN_511; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_513 = 8'hc1 == _pht2Data_T_9 ? pht_2_193 : _GEN_512; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_514 = 8'hc2 == _pht2Data_T_9 ? pht_2_194 : _GEN_513; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_515 = 8'hc3 == _pht2Data_T_9 ? pht_2_195 : _GEN_514; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_516 = 8'hc4 == _pht2Data_T_9 ? pht_2_196 : _GEN_515; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_517 = 8'hc5 == _pht2Data_T_9 ? pht_2_197 : _GEN_516; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_518 = 8'hc6 == _pht2Data_T_9 ? pht_2_198 : _GEN_517; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_519 = 8'hc7 == _pht2Data_T_9 ? pht_2_199 : _GEN_518; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_520 = 8'hc8 == _pht2Data_T_9 ? pht_2_200 : _GEN_519; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_521 = 8'hc9 == _pht2Data_T_9 ? pht_2_201 : _GEN_520; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_522 = 8'hca == _pht2Data_T_9 ? pht_2_202 : _GEN_521; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_523 = 8'hcb == _pht2Data_T_9 ? pht_2_203 : _GEN_522; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_524 = 8'hcc == _pht2Data_T_9 ? pht_2_204 : _GEN_523; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_525 = 8'hcd == _pht2Data_T_9 ? pht_2_205 : _GEN_524; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_526 = 8'hce == _pht2Data_T_9 ? pht_2_206 : _GEN_525; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_527 = 8'hcf == _pht2Data_T_9 ? pht_2_207 : _GEN_526; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_528 = 8'hd0 == _pht2Data_T_9 ? pht_2_208 : _GEN_527; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_529 = 8'hd1 == _pht2Data_T_9 ? pht_2_209 : _GEN_528; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_530 = 8'hd2 == _pht2Data_T_9 ? pht_2_210 : _GEN_529; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_531 = 8'hd3 == _pht2Data_T_9 ? pht_2_211 : _GEN_530; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_532 = 8'hd4 == _pht2Data_T_9 ? pht_2_212 : _GEN_531; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_533 = 8'hd5 == _pht2Data_T_9 ? pht_2_213 : _GEN_532; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_534 = 8'hd6 == _pht2Data_T_9 ? pht_2_214 : _GEN_533; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_535 = 8'hd7 == _pht2Data_T_9 ? pht_2_215 : _GEN_534; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_536 = 8'hd8 == _pht2Data_T_9 ? pht_2_216 : _GEN_535; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_537 = 8'hd9 == _pht2Data_T_9 ? pht_2_217 : _GEN_536; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_538 = 8'hda == _pht2Data_T_9 ? pht_2_218 : _GEN_537; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_539 = 8'hdb == _pht2Data_T_9 ? pht_2_219 : _GEN_538; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_540 = 8'hdc == _pht2Data_T_9 ? pht_2_220 : _GEN_539; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_541 = 8'hdd == _pht2Data_T_9 ? pht_2_221 : _GEN_540; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_542 = 8'hde == _pht2Data_T_9 ? pht_2_222 : _GEN_541; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_543 = 8'hdf == _pht2Data_T_9 ? pht_2_223 : _GEN_542; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_544 = 8'he0 == _pht2Data_T_9 ? pht_2_224 : _GEN_543; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_545 = 8'he1 == _pht2Data_T_9 ? pht_2_225 : _GEN_544; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_546 = 8'he2 == _pht2Data_T_9 ? pht_2_226 : _GEN_545; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_547 = 8'he3 == _pht2Data_T_9 ? pht_2_227 : _GEN_546; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_548 = 8'he4 == _pht2Data_T_9 ? pht_2_228 : _GEN_547; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_549 = 8'he5 == _pht2Data_T_9 ? pht_2_229 : _GEN_548; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_550 = 8'he6 == _pht2Data_T_9 ? pht_2_230 : _GEN_549; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_551 = 8'he7 == _pht2Data_T_9 ? pht_2_231 : _GEN_550; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_552 = 8'he8 == _pht2Data_T_9 ? pht_2_232 : _GEN_551; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_553 = 8'he9 == _pht2Data_T_9 ? pht_2_233 : _GEN_552; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_554 = 8'hea == _pht2Data_T_9 ? pht_2_234 : _GEN_553; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_555 = 8'heb == _pht2Data_T_9 ? pht_2_235 : _GEN_554; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_556 = 8'hec == _pht2Data_T_9 ? pht_2_236 : _GEN_555; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_557 = 8'hed == _pht2Data_T_9 ? pht_2_237 : _GEN_556; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_558 = 8'hee == _pht2Data_T_9 ? pht_2_238 : _GEN_557; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_559 = 8'hef == _pht2Data_T_9 ? pht_2_239 : _GEN_558; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_560 = 8'hf0 == _pht2Data_T_9 ? pht_2_240 : _GEN_559; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_561 = 8'hf1 == _pht2Data_T_9 ? pht_2_241 : _GEN_560; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_562 = 8'hf2 == _pht2Data_T_9 ? pht_2_242 : _GEN_561; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_563 = 8'hf3 == _pht2Data_T_9 ? pht_2_243 : _GEN_562; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_564 = 8'hf4 == _pht2Data_T_9 ? pht_2_244 : _GEN_563; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_565 = 8'hf5 == _pht2Data_T_9 ? pht_2_245 : _GEN_564; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_566 = 8'hf6 == _pht2Data_T_9 ? pht_2_246 : _GEN_565; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_567 = 8'hf7 == _pht2Data_T_9 ? pht_2_247 : _GEN_566; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_568 = 8'hf8 == _pht2Data_T_9 ? pht_2_248 : _GEN_567; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_569 = 8'hf9 == _pht2Data_T_9 ? pht_2_249 : _GEN_568; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_570 = 8'hfa == _pht2Data_T_9 ? pht_2_250 : _GEN_569; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_571 = 8'hfb == _pht2Data_T_9 ? pht_2_251 : _GEN_570; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_572 = 8'hfc == _pht2Data_T_9 ? pht_2_252 : _GEN_571; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_573 = 8'hfd == _pht2Data_T_9 ? pht_2_253 : _GEN_572; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_574 = 8'hfe == _pht2Data_T_9 ? pht_2_254 : _GEN_573; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_575 = 8'hff == _pht2Data_T_9 ? pht_2_255 : _GEN_574; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_577 = 8'h1 == p1Addr ? pht_1_1 : pht_1_0; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_578 = 8'h2 == p1Addr ? pht_1_2 : _GEN_577; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_579 = 8'h3 == p1Addr ? pht_1_3 : _GEN_578; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_580 = 8'h4 == p1Addr ? pht_1_4 : _GEN_579; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_581 = 8'h5 == p1Addr ? pht_1_5 : _GEN_580; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_582 = 8'h6 == p1Addr ? pht_1_6 : _GEN_581; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_583 = 8'h7 == p1Addr ? pht_1_7 : _GEN_582; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_584 = 8'h8 == p1Addr ? pht_1_8 : _GEN_583; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_585 = 8'h9 == p1Addr ? pht_1_9 : _GEN_584; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_586 = 8'ha == p1Addr ? pht_1_10 : _GEN_585; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_587 = 8'hb == p1Addr ? pht_1_11 : _GEN_586; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_588 = 8'hc == p1Addr ? pht_1_12 : _GEN_587; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_589 = 8'hd == p1Addr ? pht_1_13 : _GEN_588; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_590 = 8'he == p1Addr ? pht_1_14 : _GEN_589; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_591 = 8'hf == p1Addr ? pht_1_15 : _GEN_590; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_592 = 8'h10 == p1Addr ? pht_1_16 : _GEN_591; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_593 = 8'h11 == p1Addr ? pht_1_17 : _GEN_592; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_594 = 8'h12 == p1Addr ? pht_1_18 : _GEN_593; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_595 = 8'h13 == p1Addr ? pht_1_19 : _GEN_594; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_596 = 8'h14 == p1Addr ? pht_1_20 : _GEN_595; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_597 = 8'h15 == p1Addr ? pht_1_21 : _GEN_596; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_598 = 8'h16 == p1Addr ? pht_1_22 : _GEN_597; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_599 = 8'h17 == p1Addr ? pht_1_23 : _GEN_598; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_600 = 8'h18 == p1Addr ? pht_1_24 : _GEN_599; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_601 = 8'h19 == p1Addr ? pht_1_25 : _GEN_600; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_602 = 8'h1a == p1Addr ? pht_1_26 : _GEN_601; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_603 = 8'h1b == p1Addr ? pht_1_27 : _GEN_602; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_604 = 8'h1c == p1Addr ? pht_1_28 : _GEN_603; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_605 = 8'h1d == p1Addr ? pht_1_29 : _GEN_604; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_606 = 8'h1e == p1Addr ? pht_1_30 : _GEN_605; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_607 = 8'h1f == p1Addr ? pht_1_31 : _GEN_606; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_608 = 8'h20 == p1Addr ? pht_1_32 : _GEN_607; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_609 = 8'h21 == p1Addr ? pht_1_33 : _GEN_608; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_610 = 8'h22 == p1Addr ? pht_1_34 : _GEN_609; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_611 = 8'h23 == p1Addr ? pht_1_35 : _GEN_610; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_612 = 8'h24 == p1Addr ? pht_1_36 : _GEN_611; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_613 = 8'h25 == p1Addr ? pht_1_37 : _GEN_612; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_614 = 8'h26 == p1Addr ? pht_1_38 : _GEN_613; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_615 = 8'h27 == p1Addr ? pht_1_39 : _GEN_614; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_616 = 8'h28 == p1Addr ? pht_1_40 : _GEN_615; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_617 = 8'h29 == p1Addr ? pht_1_41 : _GEN_616; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_618 = 8'h2a == p1Addr ? pht_1_42 : _GEN_617; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_619 = 8'h2b == p1Addr ? pht_1_43 : _GEN_618; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_620 = 8'h2c == p1Addr ? pht_1_44 : _GEN_619; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_621 = 8'h2d == p1Addr ? pht_1_45 : _GEN_620; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_622 = 8'h2e == p1Addr ? pht_1_46 : _GEN_621; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_623 = 8'h2f == p1Addr ? pht_1_47 : _GEN_622; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_624 = 8'h30 == p1Addr ? pht_1_48 : _GEN_623; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_625 = 8'h31 == p1Addr ? pht_1_49 : _GEN_624; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_626 = 8'h32 == p1Addr ? pht_1_50 : _GEN_625; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_627 = 8'h33 == p1Addr ? pht_1_51 : _GEN_626; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_628 = 8'h34 == p1Addr ? pht_1_52 : _GEN_627; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_629 = 8'h35 == p1Addr ? pht_1_53 : _GEN_628; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_630 = 8'h36 == p1Addr ? pht_1_54 : _GEN_629; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_631 = 8'h37 == p1Addr ? pht_1_55 : _GEN_630; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_632 = 8'h38 == p1Addr ? pht_1_56 : _GEN_631; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_633 = 8'h39 == p1Addr ? pht_1_57 : _GEN_632; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_634 = 8'h3a == p1Addr ? pht_1_58 : _GEN_633; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_635 = 8'h3b == p1Addr ? pht_1_59 : _GEN_634; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_636 = 8'h3c == p1Addr ? pht_1_60 : _GEN_635; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_637 = 8'h3d == p1Addr ? pht_1_61 : _GEN_636; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_638 = 8'h3e == p1Addr ? pht_1_62 : _GEN_637; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_639 = 8'h3f == p1Addr ? pht_1_63 : _GEN_638; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_640 = 8'h40 == p1Addr ? pht_1_64 : _GEN_639; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_641 = 8'h41 == p1Addr ? pht_1_65 : _GEN_640; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_642 = 8'h42 == p1Addr ? pht_1_66 : _GEN_641; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_643 = 8'h43 == p1Addr ? pht_1_67 : _GEN_642; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_644 = 8'h44 == p1Addr ? pht_1_68 : _GEN_643; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_645 = 8'h45 == p1Addr ? pht_1_69 : _GEN_644; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_646 = 8'h46 == p1Addr ? pht_1_70 : _GEN_645; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_647 = 8'h47 == p1Addr ? pht_1_71 : _GEN_646; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_648 = 8'h48 == p1Addr ? pht_1_72 : _GEN_647; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_649 = 8'h49 == p1Addr ? pht_1_73 : _GEN_648; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_650 = 8'h4a == p1Addr ? pht_1_74 : _GEN_649; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_651 = 8'h4b == p1Addr ? pht_1_75 : _GEN_650; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_652 = 8'h4c == p1Addr ? pht_1_76 : _GEN_651; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_653 = 8'h4d == p1Addr ? pht_1_77 : _GEN_652; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_654 = 8'h4e == p1Addr ? pht_1_78 : _GEN_653; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_655 = 8'h4f == p1Addr ? pht_1_79 : _GEN_654; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_656 = 8'h50 == p1Addr ? pht_1_80 : _GEN_655; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_657 = 8'h51 == p1Addr ? pht_1_81 : _GEN_656; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_658 = 8'h52 == p1Addr ? pht_1_82 : _GEN_657; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_659 = 8'h53 == p1Addr ? pht_1_83 : _GEN_658; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_660 = 8'h54 == p1Addr ? pht_1_84 : _GEN_659; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_661 = 8'h55 == p1Addr ? pht_1_85 : _GEN_660; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_662 = 8'h56 == p1Addr ? pht_1_86 : _GEN_661; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_663 = 8'h57 == p1Addr ? pht_1_87 : _GEN_662; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_664 = 8'h58 == p1Addr ? pht_1_88 : _GEN_663; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_665 = 8'h59 == p1Addr ? pht_1_89 : _GEN_664; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_666 = 8'h5a == p1Addr ? pht_1_90 : _GEN_665; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_667 = 8'h5b == p1Addr ? pht_1_91 : _GEN_666; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_668 = 8'h5c == p1Addr ? pht_1_92 : _GEN_667; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_669 = 8'h5d == p1Addr ? pht_1_93 : _GEN_668; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_670 = 8'h5e == p1Addr ? pht_1_94 : _GEN_669; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_671 = 8'h5f == p1Addr ? pht_1_95 : _GEN_670; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_672 = 8'h60 == p1Addr ? pht_1_96 : _GEN_671; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_673 = 8'h61 == p1Addr ? pht_1_97 : _GEN_672; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_674 = 8'h62 == p1Addr ? pht_1_98 : _GEN_673; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_675 = 8'h63 == p1Addr ? pht_1_99 : _GEN_674; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_676 = 8'h64 == p1Addr ? pht_1_100 : _GEN_675; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_677 = 8'h65 == p1Addr ? pht_1_101 : _GEN_676; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_678 = 8'h66 == p1Addr ? pht_1_102 : _GEN_677; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_679 = 8'h67 == p1Addr ? pht_1_103 : _GEN_678; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_680 = 8'h68 == p1Addr ? pht_1_104 : _GEN_679; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_681 = 8'h69 == p1Addr ? pht_1_105 : _GEN_680; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_682 = 8'h6a == p1Addr ? pht_1_106 : _GEN_681; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_683 = 8'h6b == p1Addr ? pht_1_107 : _GEN_682; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_684 = 8'h6c == p1Addr ? pht_1_108 : _GEN_683; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_685 = 8'h6d == p1Addr ? pht_1_109 : _GEN_684; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_686 = 8'h6e == p1Addr ? pht_1_110 : _GEN_685; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_687 = 8'h6f == p1Addr ? pht_1_111 : _GEN_686; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_688 = 8'h70 == p1Addr ? pht_1_112 : _GEN_687; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_689 = 8'h71 == p1Addr ? pht_1_113 : _GEN_688; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_690 = 8'h72 == p1Addr ? pht_1_114 : _GEN_689; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_691 = 8'h73 == p1Addr ? pht_1_115 : _GEN_690; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_692 = 8'h74 == p1Addr ? pht_1_116 : _GEN_691; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_693 = 8'h75 == p1Addr ? pht_1_117 : _GEN_692; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_694 = 8'h76 == p1Addr ? pht_1_118 : _GEN_693; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_695 = 8'h77 == p1Addr ? pht_1_119 : _GEN_694; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_696 = 8'h78 == p1Addr ? pht_1_120 : _GEN_695; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_697 = 8'h79 == p1Addr ? pht_1_121 : _GEN_696; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_698 = 8'h7a == p1Addr ? pht_1_122 : _GEN_697; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_699 = 8'h7b == p1Addr ? pht_1_123 : _GEN_698; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_700 = 8'h7c == p1Addr ? pht_1_124 : _GEN_699; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_701 = 8'h7d == p1Addr ? pht_1_125 : _GEN_700; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_702 = 8'h7e == p1Addr ? pht_1_126 : _GEN_701; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_703 = 8'h7f == p1Addr ? pht_1_127 : _GEN_702; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_704 = 8'h80 == p1Addr ? pht_1_128 : _GEN_703; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_705 = 8'h81 == p1Addr ? pht_1_129 : _GEN_704; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_706 = 8'h82 == p1Addr ? pht_1_130 : _GEN_705; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_707 = 8'h83 == p1Addr ? pht_1_131 : _GEN_706; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_708 = 8'h84 == p1Addr ? pht_1_132 : _GEN_707; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_709 = 8'h85 == p1Addr ? pht_1_133 : _GEN_708; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_710 = 8'h86 == p1Addr ? pht_1_134 : _GEN_709; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_711 = 8'h87 == p1Addr ? pht_1_135 : _GEN_710; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_712 = 8'h88 == p1Addr ? pht_1_136 : _GEN_711; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_713 = 8'h89 == p1Addr ? pht_1_137 : _GEN_712; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_714 = 8'h8a == p1Addr ? pht_1_138 : _GEN_713; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_715 = 8'h8b == p1Addr ? pht_1_139 : _GEN_714; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_716 = 8'h8c == p1Addr ? pht_1_140 : _GEN_715; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_717 = 8'h8d == p1Addr ? pht_1_141 : _GEN_716; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_718 = 8'h8e == p1Addr ? pht_1_142 : _GEN_717; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_719 = 8'h8f == p1Addr ? pht_1_143 : _GEN_718; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_720 = 8'h90 == p1Addr ? pht_1_144 : _GEN_719; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_721 = 8'h91 == p1Addr ? pht_1_145 : _GEN_720; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_722 = 8'h92 == p1Addr ? pht_1_146 : _GEN_721; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_723 = 8'h93 == p1Addr ? pht_1_147 : _GEN_722; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_724 = 8'h94 == p1Addr ? pht_1_148 : _GEN_723; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_725 = 8'h95 == p1Addr ? pht_1_149 : _GEN_724; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_726 = 8'h96 == p1Addr ? pht_1_150 : _GEN_725; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_727 = 8'h97 == p1Addr ? pht_1_151 : _GEN_726; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_728 = 8'h98 == p1Addr ? pht_1_152 : _GEN_727; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_729 = 8'h99 == p1Addr ? pht_1_153 : _GEN_728; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_730 = 8'h9a == p1Addr ? pht_1_154 : _GEN_729; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_731 = 8'h9b == p1Addr ? pht_1_155 : _GEN_730; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_732 = 8'h9c == p1Addr ? pht_1_156 : _GEN_731; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_733 = 8'h9d == p1Addr ? pht_1_157 : _GEN_732; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_734 = 8'h9e == p1Addr ? pht_1_158 : _GEN_733; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_735 = 8'h9f == p1Addr ? pht_1_159 : _GEN_734; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_736 = 8'ha0 == p1Addr ? pht_1_160 : _GEN_735; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_737 = 8'ha1 == p1Addr ? pht_1_161 : _GEN_736; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_738 = 8'ha2 == p1Addr ? pht_1_162 : _GEN_737; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_739 = 8'ha3 == p1Addr ? pht_1_163 : _GEN_738; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_740 = 8'ha4 == p1Addr ? pht_1_164 : _GEN_739; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_741 = 8'ha5 == p1Addr ? pht_1_165 : _GEN_740; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_742 = 8'ha6 == p1Addr ? pht_1_166 : _GEN_741; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_743 = 8'ha7 == p1Addr ? pht_1_167 : _GEN_742; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_744 = 8'ha8 == p1Addr ? pht_1_168 : _GEN_743; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_745 = 8'ha9 == p1Addr ? pht_1_169 : _GEN_744; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_746 = 8'haa == p1Addr ? pht_1_170 : _GEN_745; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_747 = 8'hab == p1Addr ? pht_1_171 : _GEN_746; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_748 = 8'hac == p1Addr ? pht_1_172 : _GEN_747; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_749 = 8'had == p1Addr ? pht_1_173 : _GEN_748; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_750 = 8'hae == p1Addr ? pht_1_174 : _GEN_749; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_751 = 8'haf == p1Addr ? pht_1_175 : _GEN_750; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_752 = 8'hb0 == p1Addr ? pht_1_176 : _GEN_751; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_753 = 8'hb1 == p1Addr ? pht_1_177 : _GEN_752; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_754 = 8'hb2 == p1Addr ? pht_1_178 : _GEN_753; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_755 = 8'hb3 == p1Addr ? pht_1_179 : _GEN_754; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_756 = 8'hb4 == p1Addr ? pht_1_180 : _GEN_755; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_757 = 8'hb5 == p1Addr ? pht_1_181 : _GEN_756; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_758 = 8'hb6 == p1Addr ? pht_1_182 : _GEN_757; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_759 = 8'hb7 == p1Addr ? pht_1_183 : _GEN_758; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_760 = 8'hb8 == p1Addr ? pht_1_184 : _GEN_759; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_761 = 8'hb9 == p1Addr ? pht_1_185 : _GEN_760; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_762 = 8'hba == p1Addr ? pht_1_186 : _GEN_761; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_763 = 8'hbb == p1Addr ? pht_1_187 : _GEN_762; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_764 = 8'hbc == p1Addr ? pht_1_188 : _GEN_763; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_765 = 8'hbd == p1Addr ? pht_1_189 : _GEN_764; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_766 = 8'hbe == p1Addr ? pht_1_190 : _GEN_765; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_767 = 8'hbf == p1Addr ? pht_1_191 : _GEN_766; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_768 = 8'hc0 == p1Addr ? pht_1_192 : _GEN_767; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_769 = 8'hc1 == p1Addr ? pht_1_193 : _GEN_768; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_770 = 8'hc2 == p1Addr ? pht_1_194 : _GEN_769; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_771 = 8'hc3 == p1Addr ? pht_1_195 : _GEN_770; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_772 = 8'hc4 == p1Addr ? pht_1_196 : _GEN_771; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_773 = 8'hc5 == p1Addr ? pht_1_197 : _GEN_772; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_774 = 8'hc6 == p1Addr ? pht_1_198 : _GEN_773; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_775 = 8'hc7 == p1Addr ? pht_1_199 : _GEN_774; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_776 = 8'hc8 == p1Addr ? pht_1_200 : _GEN_775; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_777 = 8'hc9 == p1Addr ? pht_1_201 : _GEN_776; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_778 = 8'hca == p1Addr ? pht_1_202 : _GEN_777; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_779 = 8'hcb == p1Addr ? pht_1_203 : _GEN_778; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_780 = 8'hcc == p1Addr ? pht_1_204 : _GEN_779; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_781 = 8'hcd == p1Addr ? pht_1_205 : _GEN_780; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_782 = 8'hce == p1Addr ? pht_1_206 : _GEN_781; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_783 = 8'hcf == p1Addr ? pht_1_207 : _GEN_782; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_784 = 8'hd0 == p1Addr ? pht_1_208 : _GEN_783; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_785 = 8'hd1 == p1Addr ? pht_1_209 : _GEN_784; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_786 = 8'hd2 == p1Addr ? pht_1_210 : _GEN_785; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_787 = 8'hd3 == p1Addr ? pht_1_211 : _GEN_786; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_788 = 8'hd4 == p1Addr ? pht_1_212 : _GEN_787; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_789 = 8'hd5 == p1Addr ? pht_1_213 : _GEN_788; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_790 = 8'hd6 == p1Addr ? pht_1_214 : _GEN_789; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_791 = 8'hd7 == p1Addr ? pht_1_215 : _GEN_790; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_792 = 8'hd8 == p1Addr ? pht_1_216 : _GEN_791; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_793 = 8'hd9 == p1Addr ? pht_1_217 : _GEN_792; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_794 = 8'hda == p1Addr ? pht_1_218 : _GEN_793; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_795 = 8'hdb == p1Addr ? pht_1_219 : _GEN_794; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_796 = 8'hdc == p1Addr ? pht_1_220 : _GEN_795; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_797 = 8'hdd == p1Addr ? pht_1_221 : _GEN_796; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_798 = 8'hde == p1Addr ? pht_1_222 : _GEN_797; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_799 = 8'hdf == p1Addr ? pht_1_223 : _GEN_798; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_800 = 8'he0 == p1Addr ? pht_1_224 : _GEN_799; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_801 = 8'he1 == p1Addr ? pht_1_225 : _GEN_800; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_802 = 8'he2 == p1Addr ? pht_1_226 : _GEN_801; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_803 = 8'he3 == p1Addr ? pht_1_227 : _GEN_802; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_804 = 8'he4 == p1Addr ? pht_1_228 : _GEN_803; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_805 = 8'he5 == p1Addr ? pht_1_229 : _GEN_804; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_806 = 8'he6 == p1Addr ? pht_1_230 : _GEN_805; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_807 = 8'he7 == p1Addr ? pht_1_231 : _GEN_806; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_808 = 8'he8 == p1Addr ? pht_1_232 : _GEN_807; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_809 = 8'he9 == p1Addr ? pht_1_233 : _GEN_808; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_810 = 8'hea == p1Addr ? pht_1_234 : _GEN_809; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_811 = 8'heb == p1Addr ? pht_1_235 : _GEN_810; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_812 = 8'hec == p1Addr ? pht_1_236 : _GEN_811; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_813 = 8'hed == p1Addr ? pht_1_237 : _GEN_812; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_814 = 8'hee == p1Addr ? pht_1_238 : _GEN_813; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_815 = 8'hef == p1Addr ? pht_1_239 : _GEN_814; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_816 = 8'hf0 == p1Addr ? pht_1_240 : _GEN_815; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_817 = 8'hf1 == p1Addr ? pht_1_241 : _GEN_816; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_818 = 8'hf2 == p1Addr ? pht_1_242 : _GEN_817; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_819 = 8'hf3 == p1Addr ? pht_1_243 : _GEN_818; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_820 = 8'hf4 == p1Addr ? pht_1_244 : _GEN_819; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_821 = 8'hf5 == p1Addr ? pht_1_245 : _GEN_820; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_822 = 8'hf6 == p1Addr ? pht_1_246 : _GEN_821; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_823 = 8'hf7 == p1Addr ? pht_1_247 : _GEN_822; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_824 = 8'hf8 == p1Addr ? pht_1_248 : _GEN_823; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_825 = 8'hf9 == p1Addr ? pht_1_249 : _GEN_824; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_826 = 8'hfa == p1Addr ? pht_1_250 : _GEN_825; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_827 = 8'hfb == p1Addr ? pht_1_251 : _GEN_826; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_828 = 8'hfc == p1Addr ? pht_1_252 : _GEN_827; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_829 = 8'hfd == p1Addr ? pht_1_253 : _GEN_828; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_830 = 8'hfe == p1Addr ? pht_1_254 : _GEN_829; // @[bht.scala 60:{23,23}]
  wire [1:0] _GEN_831 = 8'hff == p1Addr ? pht_1_255 : _GEN_830; // @[bht.scala 60:{23,23}]
  wire [1:0] phtData = _GEN_319[1] ? _GEN_575 : _GEN_831; // @[bht.scala 60:23]
  reg  io_ready_REG; // @[bht.scala 64:24]
  wire [7:0] bhtWAddr_byte = io_takenPC[7:0]; // @[bht.scala 44:24]
  wire [27:0] _GEN_3341 = {{20'd0}, bhtWAddr_byte}; // @[bht.scala 45:22]
  wire [27:0] _bhtWAddr_T = 28'hce942fa ^ _GEN_3341; // @[bht.scala 45:22]
  wire [52:0] _bhtWAddr_T_1 = _bhtWAddr_T * 25'h1000193; // @[bht.scala 45:39]
  wire [7:0] bhtWAddr_byte_1 = io_takenPC[15:8]; // @[bht.scala 44:24]
  wire [52:0] _GEN_3342 = {{45'd0}, bhtWAddr_byte_1}; // @[bht.scala 45:22]
  wire [52:0] _bhtWAddr_T_2 = _bhtWAddr_T_1 ^ _GEN_3342; // @[bht.scala 45:22]
  wire [77:0] _bhtWAddr_T_3 = _bhtWAddr_T_2 * 25'h1000193; // @[bht.scala 45:39]
  wire [7:0] bhtWAddr_byte_2 = io_takenPC[23:16]; // @[bht.scala 44:24]
  wire [77:0] _GEN_3343 = {{70'd0}, bhtWAddr_byte_2}; // @[bht.scala 45:22]
  wire [77:0] _bhtWAddr_T_4 = _bhtWAddr_T_3 ^ _GEN_3343; // @[bht.scala 45:22]
  wire [102:0] _bhtWAddr_T_5 = _bhtWAddr_T_4 * 25'h1000193; // @[bht.scala 45:39]
  wire [7:0] bhtWAddr_byte_3 = io_takenPC[31:24]; // @[bht.scala 44:24]
  wire [102:0] _GEN_3344 = {{95'd0}, bhtWAddr_byte_3}; // @[bht.scala 45:22]
  wire [102:0] _bhtWAddr_T_6 = _bhtWAddr_T_5 ^ _GEN_3344; // @[bht.scala 45:22]
  wire [127:0] _bhtWAddr_T_7 = _bhtWAddr_T_6 * 25'h1000193; // @[bht.scala 45:39]
  wire [7:0] bhtWAddr = _bhtWAddr_T_7[7:0]; // @[bht.scala 49:47]
  wire [7:0] pht1WAddr = bhtWAddr ^ ghr; // @[bht.scala 50:68]
  wire [7:0] _GEN_833 = 6'h1 == bhtWAddr[5:0] ? bht_1 : bht_0; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_834 = 6'h2 == bhtWAddr[5:0] ? bht_2 : _GEN_833; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_835 = 6'h3 == bhtWAddr[5:0] ? bht_3 : _GEN_834; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_836 = 6'h4 == bhtWAddr[5:0] ? bht_4 : _GEN_835; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_837 = 6'h5 == bhtWAddr[5:0] ? bht_5 : _GEN_836; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_838 = 6'h6 == bhtWAddr[5:0] ? bht_6 : _GEN_837; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_839 = 6'h7 == bhtWAddr[5:0] ? bht_7 : _GEN_838; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_840 = 6'h8 == bhtWAddr[5:0] ? bht_8 : _GEN_839; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_841 = 6'h9 == bhtWAddr[5:0] ? bht_9 : _GEN_840; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_842 = 6'ha == bhtWAddr[5:0] ? bht_10 : _GEN_841; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_843 = 6'hb == bhtWAddr[5:0] ? bht_11 : _GEN_842; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_844 = 6'hc == bhtWAddr[5:0] ? bht_12 : _GEN_843; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_845 = 6'hd == bhtWAddr[5:0] ? bht_13 : _GEN_844; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_846 = 6'he == bhtWAddr[5:0] ? bht_14 : _GEN_845; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_847 = 6'hf == bhtWAddr[5:0] ? bht_15 : _GEN_846; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_848 = 6'h10 == bhtWAddr[5:0] ? bht_16 : _GEN_847; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_849 = 6'h11 == bhtWAddr[5:0] ? bht_17 : _GEN_848; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_850 = 6'h12 == bhtWAddr[5:0] ? bht_18 : _GEN_849; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_851 = 6'h13 == bhtWAddr[5:0] ? bht_19 : _GEN_850; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_852 = 6'h14 == bhtWAddr[5:0] ? bht_20 : _GEN_851; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_853 = 6'h15 == bhtWAddr[5:0] ? bht_21 : _GEN_852; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_854 = 6'h16 == bhtWAddr[5:0] ? bht_22 : _GEN_853; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_855 = 6'h17 == bhtWAddr[5:0] ? bht_23 : _GEN_854; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_856 = 6'h18 == bhtWAddr[5:0] ? bht_24 : _GEN_855; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_857 = 6'h19 == bhtWAddr[5:0] ? bht_25 : _GEN_856; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_858 = 6'h1a == bhtWAddr[5:0] ? bht_26 : _GEN_857; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_859 = 6'h1b == bhtWAddr[5:0] ? bht_27 : _GEN_858; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_860 = 6'h1c == bhtWAddr[5:0] ? bht_28 : _GEN_859; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_861 = 6'h1d == bhtWAddr[5:0] ? bht_29 : _GEN_860; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_862 = 6'h1e == bhtWAddr[5:0] ? bht_30 : _GEN_861; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_863 = 6'h1f == bhtWAddr[5:0] ? bht_31 : _GEN_862; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_864 = 6'h20 == bhtWAddr[5:0] ? bht_32 : _GEN_863; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_865 = 6'h21 == bhtWAddr[5:0] ? bht_33 : _GEN_864; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_866 = 6'h22 == bhtWAddr[5:0] ? bht_34 : _GEN_865; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_867 = 6'h23 == bhtWAddr[5:0] ? bht_35 : _GEN_866; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_868 = 6'h24 == bhtWAddr[5:0] ? bht_36 : _GEN_867; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_869 = 6'h25 == bhtWAddr[5:0] ? bht_37 : _GEN_868; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_870 = 6'h26 == bhtWAddr[5:0] ? bht_38 : _GEN_869; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_871 = 6'h27 == bhtWAddr[5:0] ? bht_39 : _GEN_870; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_872 = 6'h28 == bhtWAddr[5:0] ? bht_40 : _GEN_871; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_873 = 6'h29 == bhtWAddr[5:0] ? bht_41 : _GEN_872; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_874 = 6'h2a == bhtWAddr[5:0] ? bht_42 : _GEN_873; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_875 = 6'h2b == bhtWAddr[5:0] ? bht_43 : _GEN_874; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_876 = 6'h2c == bhtWAddr[5:0] ? bht_44 : _GEN_875; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_877 = 6'h2d == bhtWAddr[5:0] ? bht_45 : _GEN_876; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_878 = 6'h2e == bhtWAddr[5:0] ? bht_46 : _GEN_877; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_879 = 6'h2f == bhtWAddr[5:0] ? bht_47 : _GEN_878; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_880 = 6'h30 == bhtWAddr[5:0] ? bht_48 : _GEN_879; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_881 = 6'h31 == bhtWAddr[5:0] ? bht_49 : _GEN_880; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_882 = 6'h32 == bhtWAddr[5:0] ? bht_50 : _GEN_881; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_883 = 6'h33 == bhtWAddr[5:0] ? bht_51 : _GEN_882; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_884 = 6'h34 == bhtWAddr[5:0] ? bht_52 : _GEN_883; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_885 = 6'h35 == bhtWAddr[5:0] ? bht_53 : _GEN_884; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_886 = 6'h36 == bhtWAddr[5:0] ? bht_54 : _GEN_885; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_887 = 6'h37 == bhtWAddr[5:0] ? bht_55 : _GEN_886; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_888 = 6'h38 == bhtWAddr[5:0] ? bht_56 : _GEN_887; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_889 = 6'h39 == bhtWAddr[5:0] ? bht_57 : _GEN_888; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_890 = 6'h3a == bhtWAddr[5:0] ? bht_58 : _GEN_889; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_891 = 6'h3b == bhtWAddr[5:0] ? bht_59 : _GEN_890; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_892 = 6'h3c == bhtWAddr[5:0] ? bht_60 : _GEN_891; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_893 = 6'h3d == bhtWAddr[5:0] ? bht_61 : _GEN_892; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_894 = 6'h3e == bhtWAddr[5:0] ? bht_62 : _GEN_893; // @[bht.scala 50:{68,68}]
  wire [7:0] _GEN_895 = 6'h3f == bhtWAddr[5:0] ? bht_63 : _GEN_894; // @[bht.scala 50:{68,68}]
  wire [7:0] pht2WAddr = bhtWAddr ^ _GEN_895; // @[bht.scala 50:68]
  wire [1:0] _GEN_897 = 8'h1 == pht1WAddr ? pht_1_1 : pht_1_0; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_898 = 8'h2 == pht1WAddr ? pht_1_2 : _GEN_897; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_899 = 8'h3 == pht1WAddr ? pht_1_3 : _GEN_898; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_900 = 8'h4 == pht1WAddr ? pht_1_4 : _GEN_899; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_901 = 8'h5 == pht1WAddr ? pht_1_5 : _GEN_900; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_902 = 8'h6 == pht1WAddr ? pht_1_6 : _GEN_901; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_903 = 8'h7 == pht1WAddr ? pht_1_7 : _GEN_902; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_904 = 8'h8 == pht1WAddr ? pht_1_8 : _GEN_903; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_905 = 8'h9 == pht1WAddr ? pht_1_9 : _GEN_904; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_906 = 8'ha == pht1WAddr ? pht_1_10 : _GEN_905; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_907 = 8'hb == pht1WAddr ? pht_1_11 : _GEN_906; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_908 = 8'hc == pht1WAddr ? pht_1_12 : _GEN_907; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_909 = 8'hd == pht1WAddr ? pht_1_13 : _GEN_908; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_910 = 8'he == pht1WAddr ? pht_1_14 : _GEN_909; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_911 = 8'hf == pht1WAddr ? pht_1_15 : _GEN_910; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_912 = 8'h10 == pht1WAddr ? pht_1_16 : _GEN_911; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_913 = 8'h11 == pht1WAddr ? pht_1_17 : _GEN_912; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_914 = 8'h12 == pht1WAddr ? pht_1_18 : _GEN_913; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_915 = 8'h13 == pht1WAddr ? pht_1_19 : _GEN_914; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_916 = 8'h14 == pht1WAddr ? pht_1_20 : _GEN_915; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_917 = 8'h15 == pht1WAddr ? pht_1_21 : _GEN_916; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_918 = 8'h16 == pht1WAddr ? pht_1_22 : _GEN_917; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_919 = 8'h17 == pht1WAddr ? pht_1_23 : _GEN_918; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_920 = 8'h18 == pht1WAddr ? pht_1_24 : _GEN_919; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_921 = 8'h19 == pht1WAddr ? pht_1_25 : _GEN_920; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_922 = 8'h1a == pht1WAddr ? pht_1_26 : _GEN_921; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_923 = 8'h1b == pht1WAddr ? pht_1_27 : _GEN_922; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_924 = 8'h1c == pht1WAddr ? pht_1_28 : _GEN_923; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_925 = 8'h1d == pht1WAddr ? pht_1_29 : _GEN_924; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_926 = 8'h1e == pht1WAddr ? pht_1_30 : _GEN_925; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_927 = 8'h1f == pht1WAddr ? pht_1_31 : _GEN_926; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_928 = 8'h20 == pht1WAddr ? pht_1_32 : _GEN_927; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_929 = 8'h21 == pht1WAddr ? pht_1_33 : _GEN_928; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_930 = 8'h22 == pht1WAddr ? pht_1_34 : _GEN_929; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_931 = 8'h23 == pht1WAddr ? pht_1_35 : _GEN_930; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_932 = 8'h24 == pht1WAddr ? pht_1_36 : _GEN_931; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_933 = 8'h25 == pht1WAddr ? pht_1_37 : _GEN_932; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_934 = 8'h26 == pht1WAddr ? pht_1_38 : _GEN_933; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_935 = 8'h27 == pht1WAddr ? pht_1_39 : _GEN_934; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_936 = 8'h28 == pht1WAddr ? pht_1_40 : _GEN_935; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_937 = 8'h29 == pht1WAddr ? pht_1_41 : _GEN_936; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_938 = 8'h2a == pht1WAddr ? pht_1_42 : _GEN_937; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_939 = 8'h2b == pht1WAddr ? pht_1_43 : _GEN_938; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_940 = 8'h2c == pht1WAddr ? pht_1_44 : _GEN_939; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_941 = 8'h2d == pht1WAddr ? pht_1_45 : _GEN_940; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_942 = 8'h2e == pht1WAddr ? pht_1_46 : _GEN_941; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_943 = 8'h2f == pht1WAddr ? pht_1_47 : _GEN_942; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_944 = 8'h30 == pht1WAddr ? pht_1_48 : _GEN_943; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_945 = 8'h31 == pht1WAddr ? pht_1_49 : _GEN_944; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_946 = 8'h32 == pht1WAddr ? pht_1_50 : _GEN_945; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_947 = 8'h33 == pht1WAddr ? pht_1_51 : _GEN_946; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_948 = 8'h34 == pht1WAddr ? pht_1_52 : _GEN_947; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_949 = 8'h35 == pht1WAddr ? pht_1_53 : _GEN_948; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_950 = 8'h36 == pht1WAddr ? pht_1_54 : _GEN_949; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_951 = 8'h37 == pht1WAddr ? pht_1_55 : _GEN_950; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_952 = 8'h38 == pht1WAddr ? pht_1_56 : _GEN_951; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_953 = 8'h39 == pht1WAddr ? pht_1_57 : _GEN_952; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_954 = 8'h3a == pht1WAddr ? pht_1_58 : _GEN_953; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_955 = 8'h3b == pht1WAddr ? pht_1_59 : _GEN_954; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_956 = 8'h3c == pht1WAddr ? pht_1_60 : _GEN_955; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_957 = 8'h3d == pht1WAddr ? pht_1_61 : _GEN_956; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_958 = 8'h3e == pht1WAddr ? pht_1_62 : _GEN_957; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_959 = 8'h3f == pht1WAddr ? pht_1_63 : _GEN_958; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_960 = 8'h40 == pht1WAddr ? pht_1_64 : _GEN_959; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_961 = 8'h41 == pht1WAddr ? pht_1_65 : _GEN_960; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_962 = 8'h42 == pht1WAddr ? pht_1_66 : _GEN_961; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_963 = 8'h43 == pht1WAddr ? pht_1_67 : _GEN_962; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_964 = 8'h44 == pht1WAddr ? pht_1_68 : _GEN_963; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_965 = 8'h45 == pht1WAddr ? pht_1_69 : _GEN_964; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_966 = 8'h46 == pht1WAddr ? pht_1_70 : _GEN_965; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_967 = 8'h47 == pht1WAddr ? pht_1_71 : _GEN_966; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_968 = 8'h48 == pht1WAddr ? pht_1_72 : _GEN_967; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_969 = 8'h49 == pht1WAddr ? pht_1_73 : _GEN_968; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_970 = 8'h4a == pht1WAddr ? pht_1_74 : _GEN_969; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_971 = 8'h4b == pht1WAddr ? pht_1_75 : _GEN_970; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_972 = 8'h4c == pht1WAddr ? pht_1_76 : _GEN_971; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_973 = 8'h4d == pht1WAddr ? pht_1_77 : _GEN_972; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_974 = 8'h4e == pht1WAddr ? pht_1_78 : _GEN_973; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_975 = 8'h4f == pht1WAddr ? pht_1_79 : _GEN_974; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_976 = 8'h50 == pht1WAddr ? pht_1_80 : _GEN_975; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_977 = 8'h51 == pht1WAddr ? pht_1_81 : _GEN_976; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_978 = 8'h52 == pht1WAddr ? pht_1_82 : _GEN_977; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_979 = 8'h53 == pht1WAddr ? pht_1_83 : _GEN_978; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_980 = 8'h54 == pht1WAddr ? pht_1_84 : _GEN_979; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_981 = 8'h55 == pht1WAddr ? pht_1_85 : _GEN_980; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_982 = 8'h56 == pht1WAddr ? pht_1_86 : _GEN_981; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_983 = 8'h57 == pht1WAddr ? pht_1_87 : _GEN_982; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_984 = 8'h58 == pht1WAddr ? pht_1_88 : _GEN_983; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_985 = 8'h59 == pht1WAddr ? pht_1_89 : _GEN_984; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_986 = 8'h5a == pht1WAddr ? pht_1_90 : _GEN_985; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_987 = 8'h5b == pht1WAddr ? pht_1_91 : _GEN_986; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_988 = 8'h5c == pht1WAddr ? pht_1_92 : _GEN_987; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_989 = 8'h5d == pht1WAddr ? pht_1_93 : _GEN_988; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_990 = 8'h5e == pht1WAddr ? pht_1_94 : _GEN_989; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_991 = 8'h5f == pht1WAddr ? pht_1_95 : _GEN_990; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_992 = 8'h60 == pht1WAddr ? pht_1_96 : _GEN_991; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_993 = 8'h61 == pht1WAddr ? pht_1_97 : _GEN_992; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_994 = 8'h62 == pht1WAddr ? pht_1_98 : _GEN_993; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_995 = 8'h63 == pht1WAddr ? pht_1_99 : _GEN_994; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_996 = 8'h64 == pht1WAddr ? pht_1_100 : _GEN_995; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_997 = 8'h65 == pht1WAddr ? pht_1_101 : _GEN_996; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_998 = 8'h66 == pht1WAddr ? pht_1_102 : _GEN_997; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_999 = 8'h67 == pht1WAddr ? pht_1_103 : _GEN_998; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1000 = 8'h68 == pht1WAddr ? pht_1_104 : _GEN_999; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1001 = 8'h69 == pht1WAddr ? pht_1_105 : _GEN_1000; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1002 = 8'h6a == pht1WAddr ? pht_1_106 : _GEN_1001; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1003 = 8'h6b == pht1WAddr ? pht_1_107 : _GEN_1002; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1004 = 8'h6c == pht1WAddr ? pht_1_108 : _GEN_1003; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1005 = 8'h6d == pht1WAddr ? pht_1_109 : _GEN_1004; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1006 = 8'h6e == pht1WAddr ? pht_1_110 : _GEN_1005; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1007 = 8'h6f == pht1WAddr ? pht_1_111 : _GEN_1006; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1008 = 8'h70 == pht1WAddr ? pht_1_112 : _GEN_1007; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1009 = 8'h71 == pht1WAddr ? pht_1_113 : _GEN_1008; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1010 = 8'h72 == pht1WAddr ? pht_1_114 : _GEN_1009; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1011 = 8'h73 == pht1WAddr ? pht_1_115 : _GEN_1010; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1012 = 8'h74 == pht1WAddr ? pht_1_116 : _GEN_1011; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1013 = 8'h75 == pht1WAddr ? pht_1_117 : _GEN_1012; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1014 = 8'h76 == pht1WAddr ? pht_1_118 : _GEN_1013; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1015 = 8'h77 == pht1WAddr ? pht_1_119 : _GEN_1014; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1016 = 8'h78 == pht1WAddr ? pht_1_120 : _GEN_1015; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1017 = 8'h79 == pht1WAddr ? pht_1_121 : _GEN_1016; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1018 = 8'h7a == pht1WAddr ? pht_1_122 : _GEN_1017; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1019 = 8'h7b == pht1WAddr ? pht_1_123 : _GEN_1018; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1020 = 8'h7c == pht1WAddr ? pht_1_124 : _GEN_1019; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1021 = 8'h7d == pht1WAddr ? pht_1_125 : _GEN_1020; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1022 = 8'h7e == pht1WAddr ? pht_1_126 : _GEN_1021; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1023 = 8'h7f == pht1WAddr ? pht_1_127 : _GEN_1022; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1024 = 8'h80 == pht1WAddr ? pht_1_128 : _GEN_1023; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1025 = 8'h81 == pht1WAddr ? pht_1_129 : _GEN_1024; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1026 = 8'h82 == pht1WAddr ? pht_1_130 : _GEN_1025; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1027 = 8'h83 == pht1WAddr ? pht_1_131 : _GEN_1026; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1028 = 8'h84 == pht1WAddr ? pht_1_132 : _GEN_1027; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1029 = 8'h85 == pht1WAddr ? pht_1_133 : _GEN_1028; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1030 = 8'h86 == pht1WAddr ? pht_1_134 : _GEN_1029; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1031 = 8'h87 == pht1WAddr ? pht_1_135 : _GEN_1030; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1032 = 8'h88 == pht1WAddr ? pht_1_136 : _GEN_1031; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1033 = 8'h89 == pht1WAddr ? pht_1_137 : _GEN_1032; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1034 = 8'h8a == pht1WAddr ? pht_1_138 : _GEN_1033; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1035 = 8'h8b == pht1WAddr ? pht_1_139 : _GEN_1034; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1036 = 8'h8c == pht1WAddr ? pht_1_140 : _GEN_1035; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1037 = 8'h8d == pht1WAddr ? pht_1_141 : _GEN_1036; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1038 = 8'h8e == pht1WAddr ? pht_1_142 : _GEN_1037; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1039 = 8'h8f == pht1WAddr ? pht_1_143 : _GEN_1038; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1040 = 8'h90 == pht1WAddr ? pht_1_144 : _GEN_1039; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1041 = 8'h91 == pht1WAddr ? pht_1_145 : _GEN_1040; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1042 = 8'h92 == pht1WAddr ? pht_1_146 : _GEN_1041; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1043 = 8'h93 == pht1WAddr ? pht_1_147 : _GEN_1042; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1044 = 8'h94 == pht1WAddr ? pht_1_148 : _GEN_1043; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1045 = 8'h95 == pht1WAddr ? pht_1_149 : _GEN_1044; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1046 = 8'h96 == pht1WAddr ? pht_1_150 : _GEN_1045; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1047 = 8'h97 == pht1WAddr ? pht_1_151 : _GEN_1046; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1048 = 8'h98 == pht1WAddr ? pht_1_152 : _GEN_1047; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1049 = 8'h99 == pht1WAddr ? pht_1_153 : _GEN_1048; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1050 = 8'h9a == pht1WAddr ? pht_1_154 : _GEN_1049; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1051 = 8'h9b == pht1WAddr ? pht_1_155 : _GEN_1050; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1052 = 8'h9c == pht1WAddr ? pht_1_156 : _GEN_1051; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1053 = 8'h9d == pht1WAddr ? pht_1_157 : _GEN_1052; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1054 = 8'h9e == pht1WAddr ? pht_1_158 : _GEN_1053; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1055 = 8'h9f == pht1WAddr ? pht_1_159 : _GEN_1054; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1056 = 8'ha0 == pht1WAddr ? pht_1_160 : _GEN_1055; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1057 = 8'ha1 == pht1WAddr ? pht_1_161 : _GEN_1056; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1058 = 8'ha2 == pht1WAddr ? pht_1_162 : _GEN_1057; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1059 = 8'ha3 == pht1WAddr ? pht_1_163 : _GEN_1058; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1060 = 8'ha4 == pht1WAddr ? pht_1_164 : _GEN_1059; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1061 = 8'ha5 == pht1WAddr ? pht_1_165 : _GEN_1060; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1062 = 8'ha6 == pht1WAddr ? pht_1_166 : _GEN_1061; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1063 = 8'ha7 == pht1WAddr ? pht_1_167 : _GEN_1062; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1064 = 8'ha8 == pht1WAddr ? pht_1_168 : _GEN_1063; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1065 = 8'ha9 == pht1WAddr ? pht_1_169 : _GEN_1064; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1066 = 8'haa == pht1WAddr ? pht_1_170 : _GEN_1065; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1067 = 8'hab == pht1WAddr ? pht_1_171 : _GEN_1066; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1068 = 8'hac == pht1WAddr ? pht_1_172 : _GEN_1067; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1069 = 8'had == pht1WAddr ? pht_1_173 : _GEN_1068; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1070 = 8'hae == pht1WAddr ? pht_1_174 : _GEN_1069; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1071 = 8'haf == pht1WAddr ? pht_1_175 : _GEN_1070; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1072 = 8'hb0 == pht1WAddr ? pht_1_176 : _GEN_1071; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1073 = 8'hb1 == pht1WAddr ? pht_1_177 : _GEN_1072; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1074 = 8'hb2 == pht1WAddr ? pht_1_178 : _GEN_1073; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1075 = 8'hb3 == pht1WAddr ? pht_1_179 : _GEN_1074; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1076 = 8'hb4 == pht1WAddr ? pht_1_180 : _GEN_1075; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1077 = 8'hb5 == pht1WAddr ? pht_1_181 : _GEN_1076; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1078 = 8'hb6 == pht1WAddr ? pht_1_182 : _GEN_1077; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1079 = 8'hb7 == pht1WAddr ? pht_1_183 : _GEN_1078; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1080 = 8'hb8 == pht1WAddr ? pht_1_184 : _GEN_1079; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1081 = 8'hb9 == pht1WAddr ? pht_1_185 : _GEN_1080; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1082 = 8'hba == pht1WAddr ? pht_1_186 : _GEN_1081; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1083 = 8'hbb == pht1WAddr ? pht_1_187 : _GEN_1082; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1084 = 8'hbc == pht1WAddr ? pht_1_188 : _GEN_1083; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1085 = 8'hbd == pht1WAddr ? pht_1_189 : _GEN_1084; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1086 = 8'hbe == pht1WAddr ? pht_1_190 : _GEN_1085; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1087 = 8'hbf == pht1WAddr ? pht_1_191 : _GEN_1086; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1088 = 8'hc0 == pht1WAddr ? pht_1_192 : _GEN_1087; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1089 = 8'hc1 == pht1WAddr ? pht_1_193 : _GEN_1088; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1090 = 8'hc2 == pht1WAddr ? pht_1_194 : _GEN_1089; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1091 = 8'hc3 == pht1WAddr ? pht_1_195 : _GEN_1090; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1092 = 8'hc4 == pht1WAddr ? pht_1_196 : _GEN_1091; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1093 = 8'hc5 == pht1WAddr ? pht_1_197 : _GEN_1092; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1094 = 8'hc6 == pht1WAddr ? pht_1_198 : _GEN_1093; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1095 = 8'hc7 == pht1WAddr ? pht_1_199 : _GEN_1094; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1096 = 8'hc8 == pht1WAddr ? pht_1_200 : _GEN_1095; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1097 = 8'hc9 == pht1WAddr ? pht_1_201 : _GEN_1096; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1098 = 8'hca == pht1WAddr ? pht_1_202 : _GEN_1097; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1099 = 8'hcb == pht1WAddr ? pht_1_203 : _GEN_1098; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1100 = 8'hcc == pht1WAddr ? pht_1_204 : _GEN_1099; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1101 = 8'hcd == pht1WAddr ? pht_1_205 : _GEN_1100; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1102 = 8'hce == pht1WAddr ? pht_1_206 : _GEN_1101; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1103 = 8'hcf == pht1WAddr ? pht_1_207 : _GEN_1102; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1104 = 8'hd0 == pht1WAddr ? pht_1_208 : _GEN_1103; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1105 = 8'hd1 == pht1WAddr ? pht_1_209 : _GEN_1104; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1106 = 8'hd2 == pht1WAddr ? pht_1_210 : _GEN_1105; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1107 = 8'hd3 == pht1WAddr ? pht_1_211 : _GEN_1106; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1108 = 8'hd4 == pht1WAddr ? pht_1_212 : _GEN_1107; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1109 = 8'hd5 == pht1WAddr ? pht_1_213 : _GEN_1108; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1110 = 8'hd6 == pht1WAddr ? pht_1_214 : _GEN_1109; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1111 = 8'hd7 == pht1WAddr ? pht_1_215 : _GEN_1110; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1112 = 8'hd8 == pht1WAddr ? pht_1_216 : _GEN_1111; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1113 = 8'hd9 == pht1WAddr ? pht_1_217 : _GEN_1112; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1114 = 8'hda == pht1WAddr ? pht_1_218 : _GEN_1113; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1115 = 8'hdb == pht1WAddr ? pht_1_219 : _GEN_1114; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1116 = 8'hdc == pht1WAddr ? pht_1_220 : _GEN_1115; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1117 = 8'hdd == pht1WAddr ? pht_1_221 : _GEN_1116; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1118 = 8'hde == pht1WAddr ? pht_1_222 : _GEN_1117; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1119 = 8'hdf == pht1WAddr ? pht_1_223 : _GEN_1118; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1120 = 8'he0 == pht1WAddr ? pht_1_224 : _GEN_1119; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1121 = 8'he1 == pht1WAddr ? pht_1_225 : _GEN_1120; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1122 = 8'he2 == pht1WAddr ? pht_1_226 : _GEN_1121; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1123 = 8'he3 == pht1WAddr ? pht_1_227 : _GEN_1122; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1124 = 8'he4 == pht1WAddr ? pht_1_228 : _GEN_1123; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1125 = 8'he5 == pht1WAddr ? pht_1_229 : _GEN_1124; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1126 = 8'he6 == pht1WAddr ? pht_1_230 : _GEN_1125; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1127 = 8'he7 == pht1WAddr ? pht_1_231 : _GEN_1126; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1128 = 8'he8 == pht1WAddr ? pht_1_232 : _GEN_1127; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1129 = 8'he9 == pht1WAddr ? pht_1_233 : _GEN_1128; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1130 = 8'hea == pht1WAddr ? pht_1_234 : _GEN_1129; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1131 = 8'heb == pht1WAddr ? pht_1_235 : _GEN_1130; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1132 = 8'hec == pht1WAddr ? pht_1_236 : _GEN_1131; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1133 = 8'hed == pht1WAddr ? pht_1_237 : _GEN_1132; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1134 = 8'hee == pht1WAddr ? pht_1_238 : _GEN_1133; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1135 = 8'hef == pht1WAddr ? pht_1_239 : _GEN_1134; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1136 = 8'hf0 == pht1WAddr ? pht_1_240 : _GEN_1135; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1137 = 8'hf1 == pht1WAddr ? pht_1_241 : _GEN_1136; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1138 = 8'hf2 == pht1WAddr ? pht_1_242 : _GEN_1137; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1139 = 8'hf3 == pht1WAddr ? pht_1_243 : _GEN_1138; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1140 = 8'hf4 == pht1WAddr ? pht_1_244 : _GEN_1139; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1141 = 8'hf5 == pht1WAddr ? pht_1_245 : _GEN_1140; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1142 = 8'hf6 == pht1WAddr ? pht_1_246 : _GEN_1141; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1143 = 8'hf7 == pht1WAddr ? pht_1_247 : _GEN_1142; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1144 = 8'hf8 == pht1WAddr ? pht_1_248 : _GEN_1143; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1145 = 8'hf9 == pht1WAddr ? pht_1_249 : _GEN_1144; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1146 = 8'hfa == pht1WAddr ? pht_1_250 : _GEN_1145; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1147 = 8'hfb == pht1WAddr ? pht_1_251 : _GEN_1146; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1148 = 8'hfc == pht1WAddr ? pht_1_252 : _GEN_1147; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1149 = 8'hfd == pht1WAddr ? pht_1_253 : _GEN_1148; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1150 = 8'hfe == pht1WAddr ? pht_1_254 : _GEN_1149; // @[bht.scala 77:{26,26}]
  wire [1:0] _GEN_1151 = 8'hff == pht1WAddr ? pht_1_255 : _GEN_1150; // @[bht.scala 77:{26,26}]
  wire  p1Suc = _GEN_1151[1] == io_exTakenPre; // @[bht.scala 77:39]
  wire [1:0] _GEN_1153 = 8'h1 == pht2WAddr ? pht_2_1 : pht_2_0; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1154 = 8'h2 == pht2WAddr ? pht_2_2 : _GEN_1153; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1155 = 8'h3 == pht2WAddr ? pht_2_3 : _GEN_1154; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1156 = 8'h4 == pht2WAddr ? pht_2_4 : _GEN_1155; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1157 = 8'h5 == pht2WAddr ? pht_2_5 : _GEN_1156; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1158 = 8'h6 == pht2WAddr ? pht_2_6 : _GEN_1157; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1159 = 8'h7 == pht2WAddr ? pht_2_7 : _GEN_1158; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1160 = 8'h8 == pht2WAddr ? pht_2_8 : _GEN_1159; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1161 = 8'h9 == pht2WAddr ? pht_2_9 : _GEN_1160; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1162 = 8'ha == pht2WAddr ? pht_2_10 : _GEN_1161; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1163 = 8'hb == pht2WAddr ? pht_2_11 : _GEN_1162; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1164 = 8'hc == pht2WAddr ? pht_2_12 : _GEN_1163; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1165 = 8'hd == pht2WAddr ? pht_2_13 : _GEN_1164; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1166 = 8'he == pht2WAddr ? pht_2_14 : _GEN_1165; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1167 = 8'hf == pht2WAddr ? pht_2_15 : _GEN_1166; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1168 = 8'h10 == pht2WAddr ? pht_2_16 : _GEN_1167; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1169 = 8'h11 == pht2WAddr ? pht_2_17 : _GEN_1168; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1170 = 8'h12 == pht2WAddr ? pht_2_18 : _GEN_1169; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1171 = 8'h13 == pht2WAddr ? pht_2_19 : _GEN_1170; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1172 = 8'h14 == pht2WAddr ? pht_2_20 : _GEN_1171; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1173 = 8'h15 == pht2WAddr ? pht_2_21 : _GEN_1172; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1174 = 8'h16 == pht2WAddr ? pht_2_22 : _GEN_1173; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1175 = 8'h17 == pht2WAddr ? pht_2_23 : _GEN_1174; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1176 = 8'h18 == pht2WAddr ? pht_2_24 : _GEN_1175; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1177 = 8'h19 == pht2WAddr ? pht_2_25 : _GEN_1176; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1178 = 8'h1a == pht2WAddr ? pht_2_26 : _GEN_1177; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1179 = 8'h1b == pht2WAddr ? pht_2_27 : _GEN_1178; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1180 = 8'h1c == pht2WAddr ? pht_2_28 : _GEN_1179; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1181 = 8'h1d == pht2WAddr ? pht_2_29 : _GEN_1180; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1182 = 8'h1e == pht2WAddr ? pht_2_30 : _GEN_1181; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1183 = 8'h1f == pht2WAddr ? pht_2_31 : _GEN_1182; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1184 = 8'h20 == pht2WAddr ? pht_2_32 : _GEN_1183; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1185 = 8'h21 == pht2WAddr ? pht_2_33 : _GEN_1184; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1186 = 8'h22 == pht2WAddr ? pht_2_34 : _GEN_1185; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1187 = 8'h23 == pht2WAddr ? pht_2_35 : _GEN_1186; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1188 = 8'h24 == pht2WAddr ? pht_2_36 : _GEN_1187; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1189 = 8'h25 == pht2WAddr ? pht_2_37 : _GEN_1188; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1190 = 8'h26 == pht2WAddr ? pht_2_38 : _GEN_1189; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1191 = 8'h27 == pht2WAddr ? pht_2_39 : _GEN_1190; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1192 = 8'h28 == pht2WAddr ? pht_2_40 : _GEN_1191; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1193 = 8'h29 == pht2WAddr ? pht_2_41 : _GEN_1192; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1194 = 8'h2a == pht2WAddr ? pht_2_42 : _GEN_1193; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1195 = 8'h2b == pht2WAddr ? pht_2_43 : _GEN_1194; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1196 = 8'h2c == pht2WAddr ? pht_2_44 : _GEN_1195; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1197 = 8'h2d == pht2WAddr ? pht_2_45 : _GEN_1196; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1198 = 8'h2e == pht2WAddr ? pht_2_46 : _GEN_1197; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1199 = 8'h2f == pht2WAddr ? pht_2_47 : _GEN_1198; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1200 = 8'h30 == pht2WAddr ? pht_2_48 : _GEN_1199; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1201 = 8'h31 == pht2WAddr ? pht_2_49 : _GEN_1200; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1202 = 8'h32 == pht2WAddr ? pht_2_50 : _GEN_1201; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1203 = 8'h33 == pht2WAddr ? pht_2_51 : _GEN_1202; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1204 = 8'h34 == pht2WAddr ? pht_2_52 : _GEN_1203; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1205 = 8'h35 == pht2WAddr ? pht_2_53 : _GEN_1204; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1206 = 8'h36 == pht2WAddr ? pht_2_54 : _GEN_1205; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1207 = 8'h37 == pht2WAddr ? pht_2_55 : _GEN_1206; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1208 = 8'h38 == pht2WAddr ? pht_2_56 : _GEN_1207; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1209 = 8'h39 == pht2WAddr ? pht_2_57 : _GEN_1208; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1210 = 8'h3a == pht2WAddr ? pht_2_58 : _GEN_1209; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1211 = 8'h3b == pht2WAddr ? pht_2_59 : _GEN_1210; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1212 = 8'h3c == pht2WAddr ? pht_2_60 : _GEN_1211; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1213 = 8'h3d == pht2WAddr ? pht_2_61 : _GEN_1212; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1214 = 8'h3e == pht2WAddr ? pht_2_62 : _GEN_1213; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1215 = 8'h3f == pht2WAddr ? pht_2_63 : _GEN_1214; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1216 = 8'h40 == pht2WAddr ? pht_2_64 : _GEN_1215; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1217 = 8'h41 == pht2WAddr ? pht_2_65 : _GEN_1216; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1218 = 8'h42 == pht2WAddr ? pht_2_66 : _GEN_1217; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1219 = 8'h43 == pht2WAddr ? pht_2_67 : _GEN_1218; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1220 = 8'h44 == pht2WAddr ? pht_2_68 : _GEN_1219; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1221 = 8'h45 == pht2WAddr ? pht_2_69 : _GEN_1220; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1222 = 8'h46 == pht2WAddr ? pht_2_70 : _GEN_1221; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1223 = 8'h47 == pht2WAddr ? pht_2_71 : _GEN_1222; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1224 = 8'h48 == pht2WAddr ? pht_2_72 : _GEN_1223; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1225 = 8'h49 == pht2WAddr ? pht_2_73 : _GEN_1224; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1226 = 8'h4a == pht2WAddr ? pht_2_74 : _GEN_1225; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1227 = 8'h4b == pht2WAddr ? pht_2_75 : _GEN_1226; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1228 = 8'h4c == pht2WAddr ? pht_2_76 : _GEN_1227; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1229 = 8'h4d == pht2WAddr ? pht_2_77 : _GEN_1228; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1230 = 8'h4e == pht2WAddr ? pht_2_78 : _GEN_1229; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1231 = 8'h4f == pht2WAddr ? pht_2_79 : _GEN_1230; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1232 = 8'h50 == pht2WAddr ? pht_2_80 : _GEN_1231; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1233 = 8'h51 == pht2WAddr ? pht_2_81 : _GEN_1232; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1234 = 8'h52 == pht2WAddr ? pht_2_82 : _GEN_1233; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1235 = 8'h53 == pht2WAddr ? pht_2_83 : _GEN_1234; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1236 = 8'h54 == pht2WAddr ? pht_2_84 : _GEN_1235; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1237 = 8'h55 == pht2WAddr ? pht_2_85 : _GEN_1236; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1238 = 8'h56 == pht2WAddr ? pht_2_86 : _GEN_1237; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1239 = 8'h57 == pht2WAddr ? pht_2_87 : _GEN_1238; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1240 = 8'h58 == pht2WAddr ? pht_2_88 : _GEN_1239; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1241 = 8'h59 == pht2WAddr ? pht_2_89 : _GEN_1240; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1242 = 8'h5a == pht2WAddr ? pht_2_90 : _GEN_1241; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1243 = 8'h5b == pht2WAddr ? pht_2_91 : _GEN_1242; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1244 = 8'h5c == pht2WAddr ? pht_2_92 : _GEN_1243; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1245 = 8'h5d == pht2WAddr ? pht_2_93 : _GEN_1244; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1246 = 8'h5e == pht2WAddr ? pht_2_94 : _GEN_1245; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1247 = 8'h5f == pht2WAddr ? pht_2_95 : _GEN_1246; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1248 = 8'h60 == pht2WAddr ? pht_2_96 : _GEN_1247; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1249 = 8'h61 == pht2WAddr ? pht_2_97 : _GEN_1248; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1250 = 8'h62 == pht2WAddr ? pht_2_98 : _GEN_1249; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1251 = 8'h63 == pht2WAddr ? pht_2_99 : _GEN_1250; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1252 = 8'h64 == pht2WAddr ? pht_2_100 : _GEN_1251; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1253 = 8'h65 == pht2WAddr ? pht_2_101 : _GEN_1252; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1254 = 8'h66 == pht2WAddr ? pht_2_102 : _GEN_1253; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1255 = 8'h67 == pht2WAddr ? pht_2_103 : _GEN_1254; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1256 = 8'h68 == pht2WAddr ? pht_2_104 : _GEN_1255; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1257 = 8'h69 == pht2WAddr ? pht_2_105 : _GEN_1256; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1258 = 8'h6a == pht2WAddr ? pht_2_106 : _GEN_1257; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1259 = 8'h6b == pht2WAddr ? pht_2_107 : _GEN_1258; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1260 = 8'h6c == pht2WAddr ? pht_2_108 : _GEN_1259; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1261 = 8'h6d == pht2WAddr ? pht_2_109 : _GEN_1260; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1262 = 8'h6e == pht2WAddr ? pht_2_110 : _GEN_1261; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1263 = 8'h6f == pht2WAddr ? pht_2_111 : _GEN_1262; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1264 = 8'h70 == pht2WAddr ? pht_2_112 : _GEN_1263; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1265 = 8'h71 == pht2WAddr ? pht_2_113 : _GEN_1264; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1266 = 8'h72 == pht2WAddr ? pht_2_114 : _GEN_1265; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1267 = 8'h73 == pht2WAddr ? pht_2_115 : _GEN_1266; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1268 = 8'h74 == pht2WAddr ? pht_2_116 : _GEN_1267; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1269 = 8'h75 == pht2WAddr ? pht_2_117 : _GEN_1268; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1270 = 8'h76 == pht2WAddr ? pht_2_118 : _GEN_1269; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1271 = 8'h77 == pht2WAddr ? pht_2_119 : _GEN_1270; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1272 = 8'h78 == pht2WAddr ? pht_2_120 : _GEN_1271; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1273 = 8'h79 == pht2WAddr ? pht_2_121 : _GEN_1272; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1274 = 8'h7a == pht2WAddr ? pht_2_122 : _GEN_1273; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1275 = 8'h7b == pht2WAddr ? pht_2_123 : _GEN_1274; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1276 = 8'h7c == pht2WAddr ? pht_2_124 : _GEN_1275; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1277 = 8'h7d == pht2WAddr ? pht_2_125 : _GEN_1276; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1278 = 8'h7e == pht2WAddr ? pht_2_126 : _GEN_1277; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1279 = 8'h7f == pht2WAddr ? pht_2_127 : _GEN_1278; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1280 = 8'h80 == pht2WAddr ? pht_2_128 : _GEN_1279; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1281 = 8'h81 == pht2WAddr ? pht_2_129 : _GEN_1280; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1282 = 8'h82 == pht2WAddr ? pht_2_130 : _GEN_1281; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1283 = 8'h83 == pht2WAddr ? pht_2_131 : _GEN_1282; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1284 = 8'h84 == pht2WAddr ? pht_2_132 : _GEN_1283; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1285 = 8'h85 == pht2WAddr ? pht_2_133 : _GEN_1284; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1286 = 8'h86 == pht2WAddr ? pht_2_134 : _GEN_1285; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1287 = 8'h87 == pht2WAddr ? pht_2_135 : _GEN_1286; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1288 = 8'h88 == pht2WAddr ? pht_2_136 : _GEN_1287; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1289 = 8'h89 == pht2WAddr ? pht_2_137 : _GEN_1288; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1290 = 8'h8a == pht2WAddr ? pht_2_138 : _GEN_1289; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1291 = 8'h8b == pht2WAddr ? pht_2_139 : _GEN_1290; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1292 = 8'h8c == pht2WAddr ? pht_2_140 : _GEN_1291; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1293 = 8'h8d == pht2WAddr ? pht_2_141 : _GEN_1292; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1294 = 8'h8e == pht2WAddr ? pht_2_142 : _GEN_1293; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1295 = 8'h8f == pht2WAddr ? pht_2_143 : _GEN_1294; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1296 = 8'h90 == pht2WAddr ? pht_2_144 : _GEN_1295; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1297 = 8'h91 == pht2WAddr ? pht_2_145 : _GEN_1296; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1298 = 8'h92 == pht2WAddr ? pht_2_146 : _GEN_1297; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1299 = 8'h93 == pht2WAddr ? pht_2_147 : _GEN_1298; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1300 = 8'h94 == pht2WAddr ? pht_2_148 : _GEN_1299; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1301 = 8'h95 == pht2WAddr ? pht_2_149 : _GEN_1300; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1302 = 8'h96 == pht2WAddr ? pht_2_150 : _GEN_1301; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1303 = 8'h97 == pht2WAddr ? pht_2_151 : _GEN_1302; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1304 = 8'h98 == pht2WAddr ? pht_2_152 : _GEN_1303; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1305 = 8'h99 == pht2WAddr ? pht_2_153 : _GEN_1304; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1306 = 8'h9a == pht2WAddr ? pht_2_154 : _GEN_1305; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1307 = 8'h9b == pht2WAddr ? pht_2_155 : _GEN_1306; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1308 = 8'h9c == pht2WAddr ? pht_2_156 : _GEN_1307; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1309 = 8'h9d == pht2WAddr ? pht_2_157 : _GEN_1308; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1310 = 8'h9e == pht2WAddr ? pht_2_158 : _GEN_1309; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1311 = 8'h9f == pht2WAddr ? pht_2_159 : _GEN_1310; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1312 = 8'ha0 == pht2WAddr ? pht_2_160 : _GEN_1311; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1313 = 8'ha1 == pht2WAddr ? pht_2_161 : _GEN_1312; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1314 = 8'ha2 == pht2WAddr ? pht_2_162 : _GEN_1313; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1315 = 8'ha3 == pht2WAddr ? pht_2_163 : _GEN_1314; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1316 = 8'ha4 == pht2WAddr ? pht_2_164 : _GEN_1315; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1317 = 8'ha5 == pht2WAddr ? pht_2_165 : _GEN_1316; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1318 = 8'ha6 == pht2WAddr ? pht_2_166 : _GEN_1317; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1319 = 8'ha7 == pht2WAddr ? pht_2_167 : _GEN_1318; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1320 = 8'ha8 == pht2WAddr ? pht_2_168 : _GEN_1319; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1321 = 8'ha9 == pht2WAddr ? pht_2_169 : _GEN_1320; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1322 = 8'haa == pht2WAddr ? pht_2_170 : _GEN_1321; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1323 = 8'hab == pht2WAddr ? pht_2_171 : _GEN_1322; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1324 = 8'hac == pht2WAddr ? pht_2_172 : _GEN_1323; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1325 = 8'had == pht2WAddr ? pht_2_173 : _GEN_1324; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1326 = 8'hae == pht2WAddr ? pht_2_174 : _GEN_1325; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1327 = 8'haf == pht2WAddr ? pht_2_175 : _GEN_1326; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1328 = 8'hb0 == pht2WAddr ? pht_2_176 : _GEN_1327; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1329 = 8'hb1 == pht2WAddr ? pht_2_177 : _GEN_1328; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1330 = 8'hb2 == pht2WAddr ? pht_2_178 : _GEN_1329; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1331 = 8'hb3 == pht2WAddr ? pht_2_179 : _GEN_1330; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1332 = 8'hb4 == pht2WAddr ? pht_2_180 : _GEN_1331; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1333 = 8'hb5 == pht2WAddr ? pht_2_181 : _GEN_1332; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1334 = 8'hb6 == pht2WAddr ? pht_2_182 : _GEN_1333; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1335 = 8'hb7 == pht2WAddr ? pht_2_183 : _GEN_1334; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1336 = 8'hb8 == pht2WAddr ? pht_2_184 : _GEN_1335; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1337 = 8'hb9 == pht2WAddr ? pht_2_185 : _GEN_1336; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1338 = 8'hba == pht2WAddr ? pht_2_186 : _GEN_1337; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1339 = 8'hbb == pht2WAddr ? pht_2_187 : _GEN_1338; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1340 = 8'hbc == pht2WAddr ? pht_2_188 : _GEN_1339; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1341 = 8'hbd == pht2WAddr ? pht_2_189 : _GEN_1340; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1342 = 8'hbe == pht2WAddr ? pht_2_190 : _GEN_1341; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1343 = 8'hbf == pht2WAddr ? pht_2_191 : _GEN_1342; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1344 = 8'hc0 == pht2WAddr ? pht_2_192 : _GEN_1343; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1345 = 8'hc1 == pht2WAddr ? pht_2_193 : _GEN_1344; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1346 = 8'hc2 == pht2WAddr ? pht_2_194 : _GEN_1345; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1347 = 8'hc3 == pht2WAddr ? pht_2_195 : _GEN_1346; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1348 = 8'hc4 == pht2WAddr ? pht_2_196 : _GEN_1347; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1349 = 8'hc5 == pht2WAddr ? pht_2_197 : _GEN_1348; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1350 = 8'hc6 == pht2WAddr ? pht_2_198 : _GEN_1349; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1351 = 8'hc7 == pht2WAddr ? pht_2_199 : _GEN_1350; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1352 = 8'hc8 == pht2WAddr ? pht_2_200 : _GEN_1351; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1353 = 8'hc9 == pht2WAddr ? pht_2_201 : _GEN_1352; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1354 = 8'hca == pht2WAddr ? pht_2_202 : _GEN_1353; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1355 = 8'hcb == pht2WAddr ? pht_2_203 : _GEN_1354; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1356 = 8'hcc == pht2WAddr ? pht_2_204 : _GEN_1355; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1357 = 8'hcd == pht2WAddr ? pht_2_205 : _GEN_1356; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1358 = 8'hce == pht2WAddr ? pht_2_206 : _GEN_1357; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1359 = 8'hcf == pht2WAddr ? pht_2_207 : _GEN_1358; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1360 = 8'hd0 == pht2WAddr ? pht_2_208 : _GEN_1359; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1361 = 8'hd1 == pht2WAddr ? pht_2_209 : _GEN_1360; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1362 = 8'hd2 == pht2WAddr ? pht_2_210 : _GEN_1361; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1363 = 8'hd3 == pht2WAddr ? pht_2_211 : _GEN_1362; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1364 = 8'hd4 == pht2WAddr ? pht_2_212 : _GEN_1363; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1365 = 8'hd5 == pht2WAddr ? pht_2_213 : _GEN_1364; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1366 = 8'hd6 == pht2WAddr ? pht_2_214 : _GEN_1365; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1367 = 8'hd7 == pht2WAddr ? pht_2_215 : _GEN_1366; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1368 = 8'hd8 == pht2WAddr ? pht_2_216 : _GEN_1367; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1369 = 8'hd9 == pht2WAddr ? pht_2_217 : _GEN_1368; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1370 = 8'hda == pht2WAddr ? pht_2_218 : _GEN_1369; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1371 = 8'hdb == pht2WAddr ? pht_2_219 : _GEN_1370; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1372 = 8'hdc == pht2WAddr ? pht_2_220 : _GEN_1371; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1373 = 8'hdd == pht2WAddr ? pht_2_221 : _GEN_1372; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1374 = 8'hde == pht2WAddr ? pht_2_222 : _GEN_1373; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1375 = 8'hdf == pht2WAddr ? pht_2_223 : _GEN_1374; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1376 = 8'he0 == pht2WAddr ? pht_2_224 : _GEN_1375; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1377 = 8'he1 == pht2WAddr ? pht_2_225 : _GEN_1376; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1378 = 8'he2 == pht2WAddr ? pht_2_226 : _GEN_1377; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1379 = 8'he3 == pht2WAddr ? pht_2_227 : _GEN_1378; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1380 = 8'he4 == pht2WAddr ? pht_2_228 : _GEN_1379; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1381 = 8'he5 == pht2WAddr ? pht_2_229 : _GEN_1380; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1382 = 8'he6 == pht2WAddr ? pht_2_230 : _GEN_1381; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1383 = 8'he7 == pht2WAddr ? pht_2_231 : _GEN_1382; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1384 = 8'he8 == pht2WAddr ? pht_2_232 : _GEN_1383; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1385 = 8'he9 == pht2WAddr ? pht_2_233 : _GEN_1384; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1386 = 8'hea == pht2WAddr ? pht_2_234 : _GEN_1385; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1387 = 8'heb == pht2WAddr ? pht_2_235 : _GEN_1386; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1388 = 8'hec == pht2WAddr ? pht_2_236 : _GEN_1387; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1389 = 8'hed == pht2WAddr ? pht_2_237 : _GEN_1388; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1390 = 8'hee == pht2WAddr ? pht_2_238 : _GEN_1389; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1391 = 8'hef == pht2WAddr ? pht_2_239 : _GEN_1390; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1392 = 8'hf0 == pht2WAddr ? pht_2_240 : _GEN_1391; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1393 = 8'hf1 == pht2WAddr ? pht_2_241 : _GEN_1392; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1394 = 8'hf2 == pht2WAddr ? pht_2_242 : _GEN_1393; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1395 = 8'hf3 == pht2WAddr ? pht_2_243 : _GEN_1394; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1396 = 8'hf4 == pht2WAddr ? pht_2_244 : _GEN_1395; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1397 = 8'hf5 == pht2WAddr ? pht_2_245 : _GEN_1396; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1398 = 8'hf6 == pht2WAddr ? pht_2_246 : _GEN_1397; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1399 = 8'hf7 == pht2WAddr ? pht_2_247 : _GEN_1398; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1400 = 8'hf8 == pht2WAddr ? pht_2_248 : _GEN_1399; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1401 = 8'hf9 == pht2WAddr ? pht_2_249 : _GEN_1400; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1402 = 8'hfa == pht2WAddr ? pht_2_250 : _GEN_1401; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1403 = 8'hfb == pht2WAddr ? pht_2_251 : _GEN_1402; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1404 = 8'hfc == pht2WAddr ? pht_2_252 : _GEN_1403; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1405 = 8'hfd == pht2WAddr ? pht_2_253 : _GEN_1404; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1406 = 8'hfe == pht2WAddr ? pht_2_254 : _GEN_1405; // @[bht.scala 78:{26,26}]
  wire [1:0] _GEN_1407 = 8'hff == pht2WAddr ? pht_2_255 : _GEN_1406; // @[bht.scala 78:{26,26}]
  wire  p2Suc = _GEN_1407[1] == io_exTakenPre; // @[bht.scala 78:39]
  wire [1:0] pht0Choice = {p1Suc,p2Suc}; // @[bht.scala 79:28]
  wire  _pht_0_T = pht0Choice == 2'h1; // @[bht.scala 84:35]
  wire  _pht_0_T_3 = pht0Choice == 2'h2; // @[bht.scala 86:38]
  wire  _pht_0_T_4 = pht0Choice == 2'h2 ? 1'h0 : 1'h1; // @[bht.scala 86:26]
  wire [1:0] _pht_0_T_5 = _pht_0_T ? 2'h2 : {{1'd0}, _pht_0_T_4}; // @[bht.scala 85:23]
  wire [1:0] _pht_0_T_8 = _pht_0_T ? 2'h3 : 2'h2; // @[bht.scala 88:26]
  wire [1:0] _pht_0_T_9 = _pht_0_T_3 ? 2'h1 : _pht_0_T_8; // @[bht.scala 87:23]
  wire [1:0] _pht_0_T_11 = _pht_0_T_3 ? 2'h2 : 2'h3; // @[bht.scala 89:23]
  wire [1:0] _GEN_1409 = 8'h1 == pht1WAddr ? pht_0_1 : pht_0_0; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1410 = 8'h2 == pht1WAddr ? pht_0_2 : _GEN_1409; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1411 = 8'h3 == pht1WAddr ? pht_0_3 : _GEN_1410; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1412 = 8'h4 == pht1WAddr ? pht_0_4 : _GEN_1411; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1413 = 8'h5 == pht1WAddr ? pht_0_5 : _GEN_1412; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1414 = 8'h6 == pht1WAddr ? pht_0_6 : _GEN_1413; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1415 = 8'h7 == pht1WAddr ? pht_0_7 : _GEN_1414; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1416 = 8'h8 == pht1WAddr ? pht_0_8 : _GEN_1415; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1417 = 8'h9 == pht1WAddr ? pht_0_9 : _GEN_1416; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1418 = 8'ha == pht1WAddr ? pht_0_10 : _GEN_1417; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1419 = 8'hb == pht1WAddr ? pht_0_11 : _GEN_1418; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1420 = 8'hc == pht1WAddr ? pht_0_12 : _GEN_1419; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1421 = 8'hd == pht1WAddr ? pht_0_13 : _GEN_1420; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1422 = 8'he == pht1WAddr ? pht_0_14 : _GEN_1421; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1423 = 8'hf == pht1WAddr ? pht_0_15 : _GEN_1422; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1424 = 8'h10 == pht1WAddr ? pht_0_16 : _GEN_1423; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1425 = 8'h11 == pht1WAddr ? pht_0_17 : _GEN_1424; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1426 = 8'h12 == pht1WAddr ? pht_0_18 : _GEN_1425; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1427 = 8'h13 == pht1WAddr ? pht_0_19 : _GEN_1426; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1428 = 8'h14 == pht1WAddr ? pht_0_20 : _GEN_1427; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1429 = 8'h15 == pht1WAddr ? pht_0_21 : _GEN_1428; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1430 = 8'h16 == pht1WAddr ? pht_0_22 : _GEN_1429; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1431 = 8'h17 == pht1WAddr ? pht_0_23 : _GEN_1430; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1432 = 8'h18 == pht1WAddr ? pht_0_24 : _GEN_1431; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1433 = 8'h19 == pht1WAddr ? pht_0_25 : _GEN_1432; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1434 = 8'h1a == pht1WAddr ? pht_0_26 : _GEN_1433; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1435 = 8'h1b == pht1WAddr ? pht_0_27 : _GEN_1434; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1436 = 8'h1c == pht1WAddr ? pht_0_28 : _GEN_1435; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1437 = 8'h1d == pht1WAddr ? pht_0_29 : _GEN_1436; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1438 = 8'h1e == pht1WAddr ? pht_0_30 : _GEN_1437; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1439 = 8'h1f == pht1WAddr ? pht_0_31 : _GEN_1438; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1440 = 8'h20 == pht1WAddr ? pht_0_32 : _GEN_1439; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1441 = 8'h21 == pht1WAddr ? pht_0_33 : _GEN_1440; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1442 = 8'h22 == pht1WAddr ? pht_0_34 : _GEN_1441; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1443 = 8'h23 == pht1WAddr ? pht_0_35 : _GEN_1442; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1444 = 8'h24 == pht1WAddr ? pht_0_36 : _GEN_1443; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1445 = 8'h25 == pht1WAddr ? pht_0_37 : _GEN_1444; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1446 = 8'h26 == pht1WAddr ? pht_0_38 : _GEN_1445; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1447 = 8'h27 == pht1WAddr ? pht_0_39 : _GEN_1446; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1448 = 8'h28 == pht1WAddr ? pht_0_40 : _GEN_1447; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1449 = 8'h29 == pht1WAddr ? pht_0_41 : _GEN_1448; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1450 = 8'h2a == pht1WAddr ? pht_0_42 : _GEN_1449; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1451 = 8'h2b == pht1WAddr ? pht_0_43 : _GEN_1450; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1452 = 8'h2c == pht1WAddr ? pht_0_44 : _GEN_1451; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1453 = 8'h2d == pht1WAddr ? pht_0_45 : _GEN_1452; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1454 = 8'h2e == pht1WAddr ? pht_0_46 : _GEN_1453; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1455 = 8'h2f == pht1WAddr ? pht_0_47 : _GEN_1454; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1456 = 8'h30 == pht1WAddr ? pht_0_48 : _GEN_1455; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1457 = 8'h31 == pht1WAddr ? pht_0_49 : _GEN_1456; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1458 = 8'h32 == pht1WAddr ? pht_0_50 : _GEN_1457; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1459 = 8'h33 == pht1WAddr ? pht_0_51 : _GEN_1458; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1460 = 8'h34 == pht1WAddr ? pht_0_52 : _GEN_1459; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1461 = 8'h35 == pht1WAddr ? pht_0_53 : _GEN_1460; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1462 = 8'h36 == pht1WAddr ? pht_0_54 : _GEN_1461; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1463 = 8'h37 == pht1WAddr ? pht_0_55 : _GEN_1462; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1464 = 8'h38 == pht1WAddr ? pht_0_56 : _GEN_1463; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1465 = 8'h39 == pht1WAddr ? pht_0_57 : _GEN_1464; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1466 = 8'h3a == pht1WAddr ? pht_0_58 : _GEN_1465; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1467 = 8'h3b == pht1WAddr ? pht_0_59 : _GEN_1466; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1468 = 8'h3c == pht1WAddr ? pht_0_60 : _GEN_1467; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1469 = 8'h3d == pht1WAddr ? pht_0_61 : _GEN_1468; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1470 = 8'h3e == pht1WAddr ? pht_0_62 : _GEN_1469; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1471 = 8'h3f == pht1WAddr ? pht_0_63 : _GEN_1470; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1472 = 8'h40 == pht1WAddr ? pht_0_64 : _GEN_1471; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1473 = 8'h41 == pht1WAddr ? pht_0_65 : _GEN_1472; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1474 = 8'h42 == pht1WAddr ? pht_0_66 : _GEN_1473; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1475 = 8'h43 == pht1WAddr ? pht_0_67 : _GEN_1474; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1476 = 8'h44 == pht1WAddr ? pht_0_68 : _GEN_1475; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1477 = 8'h45 == pht1WAddr ? pht_0_69 : _GEN_1476; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1478 = 8'h46 == pht1WAddr ? pht_0_70 : _GEN_1477; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1479 = 8'h47 == pht1WAddr ? pht_0_71 : _GEN_1478; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1480 = 8'h48 == pht1WAddr ? pht_0_72 : _GEN_1479; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1481 = 8'h49 == pht1WAddr ? pht_0_73 : _GEN_1480; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1482 = 8'h4a == pht1WAddr ? pht_0_74 : _GEN_1481; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1483 = 8'h4b == pht1WAddr ? pht_0_75 : _GEN_1482; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1484 = 8'h4c == pht1WAddr ? pht_0_76 : _GEN_1483; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1485 = 8'h4d == pht1WAddr ? pht_0_77 : _GEN_1484; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1486 = 8'h4e == pht1WAddr ? pht_0_78 : _GEN_1485; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1487 = 8'h4f == pht1WAddr ? pht_0_79 : _GEN_1486; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1488 = 8'h50 == pht1WAddr ? pht_0_80 : _GEN_1487; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1489 = 8'h51 == pht1WAddr ? pht_0_81 : _GEN_1488; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1490 = 8'h52 == pht1WAddr ? pht_0_82 : _GEN_1489; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1491 = 8'h53 == pht1WAddr ? pht_0_83 : _GEN_1490; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1492 = 8'h54 == pht1WAddr ? pht_0_84 : _GEN_1491; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1493 = 8'h55 == pht1WAddr ? pht_0_85 : _GEN_1492; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1494 = 8'h56 == pht1WAddr ? pht_0_86 : _GEN_1493; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1495 = 8'h57 == pht1WAddr ? pht_0_87 : _GEN_1494; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1496 = 8'h58 == pht1WAddr ? pht_0_88 : _GEN_1495; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1497 = 8'h59 == pht1WAddr ? pht_0_89 : _GEN_1496; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1498 = 8'h5a == pht1WAddr ? pht_0_90 : _GEN_1497; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1499 = 8'h5b == pht1WAddr ? pht_0_91 : _GEN_1498; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1500 = 8'h5c == pht1WAddr ? pht_0_92 : _GEN_1499; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1501 = 8'h5d == pht1WAddr ? pht_0_93 : _GEN_1500; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1502 = 8'h5e == pht1WAddr ? pht_0_94 : _GEN_1501; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1503 = 8'h5f == pht1WAddr ? pht_0_95 : _GEN_1502; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1504 = 8'h60 == pht1WAddr ? pht_0_96 : _GEN_1503; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1505 = 8'h61 == pht1WAddr ? pht_0_97 : _GEN_1504; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1506 = 8'h62 == pht1WAddr ? pht_0_98 : _GEN_1505; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1507 = 8'h63 == pht1WAddr ? pht_0_99 : _GEN_1506; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1508 = 8'h64 == pht1WAddr ? pht_0_100 : _GEN_1507; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1509 = 8'h65 == pht1WAddr ? pht_0_101 : _GEN_1508; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1510 = 8'h66 == pht1WAddr ? pht_0_102 : _GEN_1509; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1511 = 8'h67 == pht1WAddr ? pht_0_103 : _GEN_1510; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1512 = 8'h68 == pht1WAddr ? pht_0_104 : _GEN_1511; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1513 = 8'h69 == pht1WAddr ? pht_0_105 : _GEN_1512; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1514 = 8'h6a == pht1WAddr ? pht_0_106 : _GEN_1513; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1515 = 8'h6b == pht1WAddr ? pht_0_107 : _GEN_1514; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1516 = 8'h6c == pht1WAddr ? pht_0_108 : _GEN_1515; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1517 = 8'h6d == pht1WAddr ? pht_0_109 : _GEN_1516; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1518 = 8'h6e == pht1WAddr ? pht_0_110 : _GEN_1517; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1519 = 8'h6f == pht1WAddr ? pht_0_111 : _GEN_1518; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1520 = 8'h70 == pht1WAddr ? pht_0_112 : _GEN_1519; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1521 = 8'h71 == pht1WAddr ? pht_0_113 : _GEN_1520; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1522 = 8'h72 == pht1WAddr ? pht_0_114 : _GEN_1521; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1523 = 8'h73 == pht1WAddr ? pht_0_115 : _GEN_1522; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1524 = 8'h74 == pht1WAddr ? pht_0_116 : _GEN_1523; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1525 = 8'h75 == pht1WAddr ? pht_0_117 : _GEN_1524; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1526 = 8'h76 == pht1WAddr ? pht_0_118 : _GEN_1525; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1527 = 8'h77 == pht1WAddr ? pht_0_119 : _GEN_1526; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1528 = 8'h78 == pht1WAddr ? pht_0_120 : _GEN_1527; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1529 = 8'h79 == pht1WAddr ? pht_0_121 : _GEN_1528; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1530 = 8'h7a == pht1WAddr ? pht_0_122 : _GEN_1529; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1531 = 8'h7b == pht1WAddr ? pht_0_123 : _GEN_1530; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1532 = 8'h7c == pht1WAddr ? pht_0_124 : _GEN_1531; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1533 = 8'h7d == pht1WAddr ? pht_0_125 : _GEN_1532; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1534 = 8'h7e == pht1WAddr ? pht_0_126 : _GEN_1533; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1535 = 8'h7f == pht1WAddr ? pht_0_127 : _GEN_1534; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1536 = 8'h80 == pht1WAddr ? pht_0_128 : _GEN_1535; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1537 = 8'h81 == pht1WAddr ? pht_0_129 : _GEN_1536; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1538 = 8'h82 == pht1WAddr ? pht_0_130 : _GEN_1537; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1539 = 8'h83 == pht1WAddr ? pht_0_131 : _GEN_1538; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1540 = 8'h84 == pht1WAddr ? pht_0_132 : _GEN_1539; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1541 = 8'h85 == pht1WAddr ? pht_0_133 : _GEN_1540; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1542 = 8'h86 == pht1WAddr ? pht_0_134 : _GEN_1541; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1543 = 8'h87 == pht1WAddr ? pht_0_135 : _GEN_1542; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1544 = 8'h88 == pht1WAddr ? pht_0_136 : _GEN_1543; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1545 = 8'h89 == pht1WAddr ? pht_0_137 : _GEN_1544; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1546 = 8'h8a == pht1WAddr ? pht_0_138 : _GEN_1545; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1547 = 8'h8b == pht1WAddr ? pht_0_139 : _GEN_1546; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1548 = 8'h8c == pht1WAddr ? pht_0_140 : _GEN_1547; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1549 = 8'h8d == pht1WAddr ? pht_0_141 : _GEN_1548; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1550 = 8'h8e == pht1WAddr ? pht_0_142 : _GEN_1549; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1551 = 8'h8f == pht1WAddr ? pht_0_143 : _GEN_1550; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1552 = 8'h90 == pht1WAddr ? pht_0_144 : _GEN_1551; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1553 = 8'h91 == pht1WAddr ? pht_0_145 : _GEN_1552; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1554 = 8'h92 == pht1WAddr ? pht_0_146 : _GEN_1553; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1555 = 8'h93 == pht1WAddr ? pht_0_147 : _GEN_1554; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1556 = 8'h94 == pht1WAddr ? pht_0_148 : _GEN_1555; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1557 = 8'h95 == pht1WAddr ? pht_0_149 : _GEN_1556; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1558 = 8'h96 == pht1WAddr ? pht_0_150 : _GEN_1557; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1559 = 8'h97 == pht1WAddr ? pht_0_151 : _GEN_1558; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1560 = 8'h98 == pht1WAddr ? pht_0_152 : _GEN_1559; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1561 = 8'h99 == pht1WAddr ? pht_0_153 : _GEN_1560; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1562 = 8'h9a == pht1WAddr ? pht_0_154 : _GEN_1561; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1563 = 8'h9b == pht1WAddr ? pht_0_155 : _GEN_1562; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1564 = 8'h9c == pht1WAddr ? pht_0_156 : _GEN_1563; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1565 = 8'h9d == pht1WAddr ? pht_0_157 : _GEN_1564; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1566 = 8'h9e == pht1WAddr ? pht_0_158 : _GEN_1565; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1567 = 8'h9f == pht1WAddr ? pht_0_159 : _GEN_1566; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1568 = 8'ha0 == pht1WAddr ? pht_0_160 : _GEN_1567; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1569 = 8'ha1 == pht1WAddr ? pht_0_161 : _GEN_1568; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1570 = 8'ha2 == pht1WAddr ? pht_0_162 : _GEN_1569; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1571 = 8'ha3 == pht1WAddr ? pht_0_163 : _GEN_1570; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1572 = 8'ha4 == pht1WAddr ? pht_0_164 : _GEN_1571; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1573 = 8'ha5 == pht1WAddr ? pht_0_165 : _GEN_1572; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1574 = 8'ha6 == pht1WAddr ? pht_0_166 : _GEN_1573; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1575 = 8'ha7 == pht1WAddr ? pht_0_167 : _GEN_1574; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1576 = 8'ha8 == pht1WAddr ? pht_0_168 : _GEN_1575; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1577 = 8'ha9 == pht1WAddr ? pht_0_169 : _GEN_1576; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1578 = 8'haa == pht1WAddr ? pht_0_170 : _GEN_1577; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1579 = 8'hab == pht1WAddr ? pht_0_171 : _GEN_1578; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1580 = 8'hac == pht1WAddr ? pht_0_172 : _GEN_1579; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1581 = 8'had == pht1WAddr ? pht_0_173 : _GEN_1580; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1582 = 8'hae == pht1WAddr ? pht_0_174 : _GEN_1581; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1583 = 8'haf == pht1WAddr ? pht_0_175 : _GEN_1582; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1584 = 8'hb0 == pht1WAddr ? pht_0_176 : _GEN_1583; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1585 = 8'hb1 == pht1WAddr ? pht_0_177 : _GEN_1584; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1586 = 8'hb2 == pht1WAddr ? pht_0_178 : _GEN_1585; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1587 = 8'hb3 == pht1WAddr ? pht_0_179 : _GEN_1586; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1588 = 8'hb4 == pht1WAddr ? pht_0_180 : _GEN_1587; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1589 = 8'hb5 == pht1WAddr ? pht_0_181 : _GEN_1588; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1590 = 8'hb6 == pht1WAddr ? pht_0_182 : _GEN_1589; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1591 = 8'hb7 == pht1WAddr ? pht_0_183 : _GEN_1590; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1592 = 8'hb8 == pht1WAddr ? pht_0_184 : _GEN_1591; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1593 = 8'hb9 == pht1WAddr ? pht_0_185 : _GEN_1592; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1594 = 8'hba == pht1WAddr ? pht_0_186 : _GEN_1593; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1595 = 8'hbb == pht1WAddr ? pht_0_187 : _GEN_1594; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1596 = 8'hbc == pht1WAddr ? pht_0_188 : _GEN_1595; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1597 = 8'hbd == pht1WAddr ? pht_0_189 : _GEN_1596; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1598 = 8'hbe == pht1WAddr ? pht_0_190 : _GEN_1597; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1599 = 8'hbf == pht1WAddr ? pht_0_191 : _GEN_1598; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1600 = 8'hc0 == pht1WAddr ? pht_0_192 : _GEN_1599; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1601 = 8'hc1 == pht1WAddr ? pht_0_193 : _GEN_1600; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1602 = 8'hc2 == pht1WAddr ? pht_0_194 : _GEN_1601; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1603 = 8'hc3 == pht1WAddr ? pht_0_195 : _GEN_1602; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1604 = 8'hc4 == pht1WAddr ? pht_0_196 : _GEN_1603; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1605 = 8'hc5 == pht1WAddr ? pht_0_197 : _GEN_1604; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1606 = 8'hc6 == pht1WAddr ? pht_0_198 : _GEN_1605; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1607 = 8'hc7 == pht1WAddr ? pht_0_199 : _GEN_1606; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1608 = 8'hc8 == pht1WAddr ? pht_0_200 : _GEN_1607; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1609 = 8'hc9 == pht1WAddr ? pht_0_201 : _GEN_1608; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1610 = 8'hca == pht1WAddr ? pht_0_202 : _GEN_1609; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1611 = 8'hcb == pht1WAddr ? pht_0_203 : _GEN_1610; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1612 = 8'hcc == pht1WAddr ? pht_0_204 : _GEN_1611; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1613 = 8'hcd == pht1WAddr ? pht_0_205 : _GEN_1612; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1614 = 8'hce == pht1WAddr ? pht_0_206 : _GEN_1613; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1615 = 8'hcf == pht1WAddr ? pht_0_207 : _GEN_1614; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1616 = 8'hd0 == pht1WAddr ? pht_0_208 : _GEN_1615; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1617 = 8'hd1 == pht1WAddr ? pht_0_209 : _GEN_1616; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1618 = 8'hd2 == pht1WAddr ? pht_0_210 : _GEN_1617; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1619 = 8'hd3 == pht1WAddr ? pht_0_211 : _GEN_1618; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1620 = 8'hd4 == pht1WAddr ? pht_0_212 : _GEN_1619; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1621 = 8'hd5 == pht1WAddr ? pht_0_213 : _GEN_1620; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1622 = 8'hd6 == pht1WAddr ? pht_0_214 : _GEN_1621; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1623 = 8'hd7 == pht1WAddr ? pht_0_215 : _GEN_1622; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1624 = 8'hd8 == pht1WAddr ? pht_0_216 : _GEN_1623; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1625 = 8'hd9 == pht1WAddr ? pht_0_217 : _GEN_1624; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1626 = 8'hda == pht1WAddr ? pht_0_218 : _GEN_1625; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1627 = 8'hdb == pht1WAddr ? pht_0_219 : _GEN_1626; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1628 = 8'hdc == pht1WAddr ? pht_0_220 : _GEN_1627; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1629 = 8'hdd == pht1WAddr ? pht_0_221 : _GEN_1628; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1630 = 8'hde == pht1WAddr ? pht_0_222 : _GEN_1629; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1631 = 8'hdf == pht1WAddr ? pht_0_223 : _GEN_1630; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1632 = 8'he0 == pht1WAddr ? pht_0_224 : _GEN_1631; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1633 = 8'he1 == pht1WAddr ? pht_0_225 : _GEN_1632; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1634 = 8'he2 == pht1WAddr ? pht_0_226 : _GEN_1633; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1635 = 8'he3 == pht1WAddr ? pht_0_227 : _GEN_1634; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1636 = 8'he4 == pht1WAddr ? pht_0_228 : _GEN_1635; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1637 = 8'he5 == pht1WAddr ? pht_0_229 : _GEN_1636; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1638 = 8'he6 == pht1WAddr ? pht_0_230 : _GEN_1637; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1639 = 8'he7 == pht1WAddr ? pht_0_231 : _GEN_1638; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1640 = 8'he8 == pht1WAddr ? pht_0_232 : _GEN_1639; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1641 = 8'he9 == pht1WAddr ? pht_0_233 : _GEN_1640; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1642 = 8'hea == pht1WAddr ? pht_0_234 : _GEN_1641; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1643 = 8'heb == pht1WAddr ? pht_0_235 : _GEN_1642; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1644 = 8'hec == pht1WAddr ? pht_0_236 : _GEN_1643; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1645 = 8'hed == pht1WAddr ? pht_0_237 : _GEN_1644; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1646 = 8'hee == pht1WAddr ? pht_0_238 : _GEN_1645; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1647 = 8'hef == pht1WAddr ? pht_0_239 : _GEN_1646; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1648 = 8'hf0 == pht1WAddr ? pht_0_240 : _GEN_1647; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1649 = 8'hf1 == pht1WAddr ? pht_0_241 : _GEN_1648; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1650 = 8'hf2 == pht1WAddr ? pht_0_242 : _GEN_1649; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1651 = 8'hf3 == pht1WAddr ? pht_0_243 : _GEN_1650; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1652 = 8'hf4 == pht1WAddr ? pht_0_244 : _GEN_1651; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1653 = 8'hf5 == pht1WAddr ? pht_0_245 : _GEN_1652; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1654 = 8'hf6 == pht1WAddr ? pht_0_246 : _GEN_1653; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1655 = 8'hf7 == pht1WAddr ? pht_0_247 : _GEN_1654; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1656 = 8'hf8 == pht1WAddr ? pht_0_248 : _GEN_1655; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1657 = 8'hf9 == pht1WAddr ? pht_0_249 : _GEN_1656; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1658 = 8'hfa == pht1WAddr ? pht_0_250 : _GEN_1657; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1659 = 8'hfb == pht1WAddr ? pht_0_251 : _GEN_1658; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1660 = 8'hfc == pht1WAddr ? pht_0_252 : _GEN_1659; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1661 = 8'hfd == pht1WAddr ? pht_0_253 : _GEN_1660; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1662 = 8'hfe == pht1WAddr ? pht_0_254 : _GEN_1661; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1663 = 8'hff == pht1WAddr ? pht_0_255 : _GEN_1662; // @[Mux.scala 81:{61,61}]
  wire [1:0] _pht_0_T_13 = 2'h1 == _GEN_1663 ? _pht_0_T_5 : {{1'd0}, _pht_0_T}; // @[Mux.scala 81:58]
  wire [1:0] _pht_0_T_15 = 2'h2 == _GEN_1663 ? _pht_0_T_9 : _pht_0_T_13; // @[Mux.scala 81:58]
  wire [1:0] _pht_1_T_1 = io_takenMiss ? 2'h2 : 2'h0; // @[bht.scala 95:23]
  wire [1:0] _pht_1_T_2 = io_takenMiss ? 2'h1 : 2'h3; // @[bht.scala 96:23]
  wire [1:0] _pht_1_T_3 = io_takenMiss ? 2'h2 : 2'h3; // @[bht.scala 97:23]
  wire [1:0] _pht_1_T_5 = 2'h1 == _GEN_1151 ? _pht_1_T_1 : {{1'd0}, io_takenMiss}; // @[Mux.scala 81:58]
  wire [1:0] _pht_1_T_7 = 2'h2 == _GEN_1151 ? _pht_1_T_2 : _pht_1_T_5; // @[Mux.scala 81:58]
  wire [1:0] _pht_2_T_5 = 2'h1 == _GEN_1407 ? _pht_1_T_1 : {{1'd0}, io_takenMiss}; // @[Mux.scala 81:58]
  wire [1:0] _pht_2_T_7 = 2'h2 == _GEN_1407 ? _pht_1_T_2 : _pht_2_T_5; // @[Mux.scala 81:58]
  wire [7:0] _bht_T_1 = {_GEN_895[6:0],io_exTakenPre}; // @[bht.scala 110:49]
  wire [7:0] _ghr_T_1 = {ghr[6:0],io_exTakenPre}; // @[bht.scala 111:33]
  assign io_takenPre = io_valid & phtData[1]; // @[bht.scala 63:23]
  assign io_ready = io_ready_REG; // @[bht.scala 64:14]
  always @(posedge clock) begin
    if (reset) begin // @[bht.scala 51:22]
      ghr <= 8'h0; // @[bht.scala 51:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      ghr <= _ghr_T_1; // @[bht.scala 111:11]
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_0 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h0 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_0 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_1 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h1 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_1 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_2 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h2 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_2 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_3 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h3 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_3 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_4 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h4 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_4 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_5 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h5 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_5 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_6 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h6 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_6 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_7 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h7 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_7 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_8 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h8 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_8 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_9 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h9 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_9 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_10 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'ha == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_10 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_11 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'hb == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_11 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_12 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'hc == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_12 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_13 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'hd == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_13 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_14 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'he == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_14 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_15 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'hf == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_15 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_16 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h10 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_16 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_17 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h11 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_17 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_18 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h12 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_18 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_19 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h13 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_19 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_20 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h14 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_20 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_21 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h15 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_21 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_22 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h16 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_22 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_23 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h17 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_23 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_24 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h18 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_24 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_25 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h19 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_25 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_26 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h1a == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_26 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_27 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h1b == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_27 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_28 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h1c == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_28 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_29 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h1d == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_29 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_30 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h1e == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_30 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_31 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h1f == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_31 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_32 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h20 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_32 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_33 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h21 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_33 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_34 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h22 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_34 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_35 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h23 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_35 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_36 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h24 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_36 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_37 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h25 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_37 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_38 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h26 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_38 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_39 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h27 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_39 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_40 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h28 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_40 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_41 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h29 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_41 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_42 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h2a == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_42 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_43 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h2b == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_43 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_44 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h2c == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_44 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_45 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h2d == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_45 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_46 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h2e == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_46 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_47 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h2f == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_47 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_48 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h30 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_48 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_49 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h31 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_49 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_50 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h32 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_50 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_51 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h33 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_51 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_52 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h34 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_52 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_53 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h35 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_53 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_54 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h36 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_54 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_55 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h37 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_55 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_56 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h38 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_56 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_57 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h39 == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_57 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_58 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h3a == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_58 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_59 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h3b == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_59 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_60 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h3c == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_60 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_61 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h3d == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_61 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_62 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h3e == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_62 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 52:22]
      bht_63 <= 8'h0; // @[bht.scala 52:22]
    end else if (io_takenValid) begin // @[bht.scala 109:25]
      if (6'h3f == bhtWAddr[5:0]) begin // @[bht.scala 110:21]
        bht_63 <= _bht_T_1; // @[bht.scala 110:21]
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_0 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h0 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_0 <= _pht_0_T_11;
        end else begin
          pht_0_0 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_1 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h1 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_1 <= _pht_0_T_11;
        end else begin
          pht_0_1 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_2 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h2 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_2 <= _pht_0_T_11;
        end else begin
          pht_0_2 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_3 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h3 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_3 <= _pht_0_T_11;
        end else begin
          pht_0_3 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_4 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h4 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_4 <= _pht_0_T_11;
        end else begin
          pht_0_4 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_5 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h5 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_5 <= _pht_0_T_11;
        end else begin
          pht_0_5 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_6 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h6 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_6 <= _pht_0_T_11;
        end else begin
          pht_0_6 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_7 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h7 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_7 <= _pht_0_T_11;
        end else begin
          pht_0_7 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_8 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h8 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_8 <= _pht_0_T_11;
        end else begin
          pht_0_8 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_9 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h9 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_9 <= _pht_0_T_11;
        end else begin
          pht_0_9 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_10 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_10 <= _pht_0_T_11;
        end else begin
          pht_0_10 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_11 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_11 <= _pht_0_T_11;
        end else begin
          pht_0_11 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_12 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_12 <= _pht_0_T_11;
        end else begin
          pht_0_12 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_13 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_13 <= _pht_0_T_11;
        end else begin
          pht_0_13 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_14 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_14 <= _pht_0_T_11;
        end else begin
          pht_0_14 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_15 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_15 <= _pht_0_T_11;
        end else begin
          pht_0_15 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_16 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h10 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_16 <= _pht_0_T_11;
        end else begin
          pht_0_16 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_17 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h11 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_17 <= _pht_0_T_11;
        end else begin
          pht_0_17 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_18 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h12 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_18 <= _pht_0_T_11;
        end else begin
          pht_0_18 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_19 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h13 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_19 <= _pht_0_T_11;
        end else begin
          pht_0_19 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_20 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h14 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_20 <= _pht_0_T_11;
        end else begin
          pht_0_20 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_21 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h15 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_21 <= _pht_0_T_11;
        end else begin
          pht_0_21 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_22 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h16 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_22 <= _pht_0_T_11;
        end else begin
          pht_0_22 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_23 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h17 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_23 <= _pht_0_T_11;
        end else begin
          pht_0_23 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_24 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h18 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_24 <= _pht_0_T_11;
        end else begin
          pht_0_24 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_25 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h19 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_25 <= _pht_0_T_11;
        end else begin
          pht_0_25 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_26 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h1a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_26 <= _pht_0_T_11;
        end else begin
          pht_0_26 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_27 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h1b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_27 <= _pht_0_T_11;
        end else begin
          pht_0_27 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_28 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h1c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_28 <= _pht_0_T_11;
        end else begin
          pht_0_28 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_29 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h1d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_29 <= _pht_0_T_11;
        end else begin
          pht_0_29 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_30 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h1e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_30 <= _pht_0_T_11;
        end else begin
          pht_0_30 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_31 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h1f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_31 <= _pht_0_T_11;
        end else begin
          pht_0_31 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_32 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h20 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_32 <= _pht_0_T_11;
        end else begin
          pht_0_32 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_33 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h21 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_33 <= _pht_0_T_11;
        end else begin
          pht_0_33 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_34 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h22 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_34 <= _pht_0_T_11;
        end else begin
          pht_0_34 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_35 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h23 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_35 <= _pht_0_T_11;
        end else begin
          pht_0_35 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_36 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h24 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_36 <= _pht_0_T_11;
        end else begin
          pht_0_36 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_37 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h25 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_37 <= _pht_0_T_11;
        end else begin
          pht_0_37 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_38 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h26 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_38 <= _pht_0_T_11;
        end else begin
          pht_0_38 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_39 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h27 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_39 <= _pht_0_T_11;
        end else begin
          pht_0_39 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_40 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h28 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_40 <= _pht_0_T_11;
        end else begin
          pht_0_40 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_41 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h29 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_41 <= _pht_0_T_11;
        end else begin
          pht_0_41 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_42 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h2a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_42 <= _pht_0_T_11;
        end else begin
          pht_0_42 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_43 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h2b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_43 <= _pht_0_T_11;
        end else begin
          pht_0_43 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_44 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h2c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_44 <= _pht_0_T_11;
        end else begin
          pht_0_44 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_45 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h2d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_45 <= _pht_0_T_11;
        end else begin
          pht_0_45 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_46 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h2e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_46 <= _pht_0_T_11;
        end else begin
          pht_0_46 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_47 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h2f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_47 <= _pht_0_T_11;
        end else begin
          pht_0_47 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_48 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h30 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_48 <= _pht_0_T_11;
        end else begin
          pht_0_48 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_49 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h31 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_49 <= _pht_0_T_11;
        end else begin
          pht_0_49 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_50 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h32 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_50 <= _pht_0_T_11;
        end else begin
          pht_0_50 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_51 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h33 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_51 <= _pht_0_T_11;
        end else begin
          pht_0_51 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_52 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h34 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_52 <= _pht_0_T_11;
        end else begin
          pht_0_52 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_53 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h35 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_53 <= _pht_0_T_11;
        end else begin
          pht_0_53 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_54 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h36 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_54 <= _pht_0_T_11;
        end else begin
          pht_0_54 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_55 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h37 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_55 <= _pht_0_T_11;
        end else begin
          pht_0_55 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_56 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h38 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_56 <= _pht_0_T_11;
        end else begin
          pht_0_56 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_57 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h39 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_57 <= _pht_0_T_11;
        end else begin
          pht_0_57 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_58 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h3a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_58 <= _pht_0_T_11;
        end else begin
          pht_0_58 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_59 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h3b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_59 <= _pht_0_T_11;
        end else begin
          pht_0_59 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_60 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h3c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_60 <= _pht_0_T_11;
        end else begin
          pht_0_60 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_61 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h3d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_61 <= _pht_0_T_11;
        end else begin
          pht_0_61 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_62 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h3e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_62 <= _pht_0_T_11;
        end else begin
          pht_0_62 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_63 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h3f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_63 <= _pht_0_T_11;
        end else begin
          pht_0_63 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_64 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h40 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_64 <= _pht_0_T_11;
        end else begin
          pht_0_64 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_65 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h41 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_65 <= _pht_0_T_11;
        end else begin
          pht_0_65 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_66 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h42 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_66 <= _pht_0_T_11;
        end else begin
          pht_0_66 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_67 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h43 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_67 <= _pht_0_T_11;
        end else begin
          pht_0_67 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_68 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h44 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_68 <= _pht_0_T_11;
        end else begin
          pht_0_68 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_69 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h45 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_69 <= _pht_0_T_11;
        end else begin
          pht_0_69 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_70 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h46 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_70 <= _pht_0_T_11;
        end else begin
          pht_0_70 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_71 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h47 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_71 <= _pht_0_T_11;
        end else begin
          pht_0_71 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_72 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h48 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_72 <= _pht_0_T_11;
        end else begin
          pht_0_72 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_73 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h49 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_73 <= _pht_0_T_11;
        end else begin
          pht_0_73 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_74 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h4a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_74 <= _pht_0_T_11;
        end else begin
          pht_0_74 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_75 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h4b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_75 <= _pht_0_T_11;
        end else begin
          pht_0_75 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_76 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h4c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_76 <= _pht_0_T_11;
        end else begin
          pht_0_76 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_77 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h4d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_77 <= _pht_0_T_11;
        end else begin
          pht_0_77 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_78 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h4e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_78 <= _pht_0_T_11;
        end else begin
          pht_0_78 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_79 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h4f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_79 <= _pht_0_T_11;
        end else begin
          pht_0_79 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_80 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h50 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_80 <= _pht_0_T_11;
        end else begin
          pht_0_80 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_81 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h51 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_81 <= _pht_0_T_11;
        end else begin
          pht_0_81 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_82 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h52 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_82 <= _pht_0_T_11;
        end else begin
          pht_0_82 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_83 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h53 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_83 <= _pht_0_T_11;
        end else begin
          pht_0_83 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_84 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h54 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_84 <= _pht_0_T_11;
        end else begin
          pht_0_84 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_85 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h55 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_85 <= _pht_0_T_11;
        end else begin
          pht_0_85 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_86 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h56 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_86 <= _pht_0_T_11;
        end else begin
          pht_0_86 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_87 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h57 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_87 <= _pht_0_T_11;
        end else begin
          pht_0_87 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_88 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h58 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_88 <= _pht_0_T_11;
        end else begin
          pht_0_88 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_89 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h59 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_89 <= _pht_0_T_11;
        end else begin
          pht_0_89 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_90 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h5a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_90 <= _pht_0_T_11;
        end else begin
          pht_0_90 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_91 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h5b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_91 <= _pht_0_T_11;
        end else begin
          pht_0_91 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_92 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h5c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_92 <= _pht_0_T_11;
        end else begin
          pht_0_92 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_93 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h5d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_93 <= _pht_0_T_11;
        end else begin
          pht_0_93 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_94 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h5e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_94 <= _pht_0_T_11;
        end else begin
          pht_0_94 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_95 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h5f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_95 <= _pht_0_T_11;
        end else begin
          pht_0_95 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_96 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h60 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_96 <= _pht_0_T_11;
        end else begin
          pht_0_96 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_97 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h61 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_97 <= _pht_0_T_11;
        end else begin
          pht_0_97 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_98 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h62 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_98 <= _pht_0_T_11;
        end else begin
          pht_0_98 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_99 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h63 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_99 <= _pht_0_T_11;
        end else begin
          pht_0_99 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_100 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h64 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_100 <= _pht_0_T_11;
        end else begin
          pht_0_100 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_101 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h65 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_101 <= _pht_0_T_11;
        end else begin
          pht_0_101 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_102 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h66 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_102 <= _pht_0_T_11;
        end else begin
          pht_0_102 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_103 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h67 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_103 <= _pht_0_T_11;
        end else begin
          pht_0_103 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_104 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h68 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_104 <= _pht_0_T_11;
        end else begin
          pht_0_104 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_105 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h69 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_105 <= _pht_0_T_11;
        end else begin
          pht_0_105 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_106 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h6a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_106 <= _pht_0_T_11;
        end else begin
          pht_0_106 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_107 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h6b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_107 <= _pht_0_T_11;
        end else begin
          pht_0_107 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_108 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h6c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_108 <= _pht_0_T_11;
        end else begin
          pht_0_108 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_109 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h6d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_109 <= _pht_0_T_11;
        end else begin
          pht_0_109 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_110 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h6e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_110 <= _pht_0_T_11;
        end else begin
          pht_0_110 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_111 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h6f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_111 <= _pht_0_T_11;
        end else begin
          pht_0_111 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_112 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h70 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_112 <= _pht_0_T_11;
        end else begin
          pht_0_112 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_113 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h71 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_113 <= _pht_0_T_11;
        end else begin
          pht_0_113 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_114 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h72 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_114 <= _pht_0_T_11;
        end else begin
          pht_0_114 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_115 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h73 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_115 <= _pht_0_T_11;
        end else begin
          pht_0_115 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_116 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h74 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_116 <= _pht_0_T_11;
        end else begin
          pht_0_116 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_117 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h75 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_117 <= _pht_0_T_11;
        end else begin
          pht_0_117 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_118 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h76 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_118 <= _pht_0_T_11;
        end else begin
          pht_0_118 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_119 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h77 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_119 <= _pht_0_T_11;
        end else begin
          pht_0_119 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_120 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h78 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_120 <= _pht_0_T_11;
        end else begin
          pht_0_120 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_121 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h79 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_121 <= _pht_0_T_11;
        end else begin
          pht_0_121 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_122 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h7a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_122 <= _pht_0_T_11;
        end else begin
          pht_0_122 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_123 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h7b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_123 <= _pht_0_T_11;
        end else begin
          pht_0_123 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_124 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h7c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_124 <= _pht_0_T_11;
        end else begin
          pht_0_124 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_125 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h7d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_125 <= _pht_0_T_11;
        end else begin
          pht_0_125 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_126 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h7e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_126 <= _pht_0_T_11;
        end else begin
          pht_0_126 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_127 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h7f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_127 <= _pht_0_T_11;
        end else begin
          pht_0_127 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_128 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h80 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_128 <= _pht_0_T_11;
        end else begin
          pht_0_128 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_129 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h81 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_129 <= _pht_0_T_11;
        end else begin
          pht_0_129 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_130 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h82 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_130 <= _pht_0_T_11;
        end else begin
          pht_0_130 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_131 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h83 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_131 <= _pht_0_T_11;
        end else begin
          pht_0_131 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_132 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h84 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_132 <= _pht_0_T_11;
        end else begin
          pht_0_132 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_133 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h85 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_133 <= _pht_0_T_11;
        end else begin
          pht_0_133 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_134 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h86 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_134 <= _pht_0_T_11;
        end else begin
          pht_0_134 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_135 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h87 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_135 <= _pht_0_T_11;
        end else begin
          pht_0_135 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_136 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h88 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_136 <= _pht_0_T_11;
        end else begin
          pht_0_136 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_137 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h89 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_137 <= _pht_0_T_11;
        end else begin
          pht_0_137 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_138 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h8a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_138 <= _pht_0_T_11;
        end else begin
          pht_0_138 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_139 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h8b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_139 <= _pht_0_T_11;
        end else begin
          pht_0_139 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_140 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h8c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_140 <= _pht_0_T_11;
        end else begin
          pht_0_140 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_141 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h8d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_141 <= _pht_0_T_11;
        end else begin
          pht_0_141 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_142 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h8e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_142 <= _pht_0_T_11;
        end else begin
          pht_0_142 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_143 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h8f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_143 <= _pht_0_T_11;
        end else begin
          pht_0_143 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_144 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h90 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_144 <= _pht_0_T_11;
        end else begin
          pht_0_144 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_145 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h91 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_145 <= _pht_0_T_11;
        end else begin
          pht_0_145 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_146 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h92 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_146 <= _pht_0_T_11;
        end else begin
          pht_0_146 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_147 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h93 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_147 <= _pht_0_T_11;
        end else begin
          pht_0_147 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_148 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h94 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_148 <= _pht_0_T_11;
        end else begin
          pht_0_148 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_149 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h95 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_149 <= _pht_0_T_11;
        end else begin
          pht_0_149 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_150 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h96 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_150 <= _pht_0_T_11;
        end else begin
          pht_0_150 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_151 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h97 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_151 <= _pht_0_T_11;
        end else begin
          pht_0_151 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_152 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h98 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_152 <= _pht_0_T_11;
        end else begin
          pht_0_152 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_153 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h99 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_153 <= _pht_0_T_11;
        end else begin
          pht_0_153 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_154 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h9a == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_154 <= _pht_0_T_11;
        end else begin
          pht_0_154 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_155 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h9b == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_155 <= _pht_0_T_11;
        end else begin
          pht_0_155 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_156 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h9c == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_156 <= _pht_0_T_11;
        end else begin
          pht_0_156 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_157 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h9d == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_157 <= _pht_0_T_11;
        end else begin
          pht_0_157 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_158 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h9e == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_158 <= _pht_0_T_11;
        end else begin
          pht_0_158 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_159 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'h9f == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_159 <= _pht_0_T_11;
        end else begin
          pht_0_159 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_160 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha0 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_160 <= _pht_0_T_11;
        end else begin
          pht_0_160 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_161 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha1 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_161 <= _pht_0_T_11;
        end else begin
          pht_0_161 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_162 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha2 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_162 <= _pht_0_T_11;
        end else begin
          pht_0_162 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_163 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha3 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_163 <= _pht_0_T_11;
        end else begin
          pht_0_163 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_164 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha4 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_164 <= _pht_0_T_11;
        end else begin
          pht_0_164 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_165 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha5 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_165 <= _pht_0_T_11;
        end else begin
          pht_0_165 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_166 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha6 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_166 <= _pht_0_T_11;
        end else begin
          pht_0_166 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_167 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha7 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_167 <= _pht_0_T_11;
        end else begin
          pht_0_167 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_168 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha8 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_168 <= _pht_0_T_11;
        end else begin
          pht_0_168 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_169 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'ha9 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_169 <= _pht_0_T_11;
        end else begin
          pht_0_169 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_170 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'haa == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_170 <= _pht_0_T_11;
        end else begin
          pht_0_170 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_171 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hab == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_171 <= _pht_0_T_11;
        end else begin
          pht_0_171 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_172 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hac == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_172 <= _pht_0_T_11;
        end else begin
          pht_0_172 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_173 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'had == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_173 <= _pht_0_T_11;
        end else begin
          pht_0_173 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_174 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hae == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_174 <= _pht_0_T_11;
        end else begin
          pht_0_174 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_175 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'haf == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_175 <= _pht_0_T_11;
        end else begin
          pht_0_175 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_176 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb0 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_176 <= _pht_0_T_11;
        end else begin
          pht_0_176 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_177 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb1 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_177 <= _pht_0_T_11;
        end else begin
          pht_0_177 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_178 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb2 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_178 <= _pht_0_T_11;
        end else begin
          pht_0_178 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_179 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb3 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_179 <= _pht_0_T_11;
        end else begin
          pht_0_179 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_180 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb4 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_180 <= _pht_0_T_11;
        end else begin
          pht_0_180 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_181 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb5 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_181 <= _pht_0_T_11;
        end else begin
          pht_0_181 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_182 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb6 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_182 <= _pht_0_T_11;
        end else begin
          pht_0_182 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_183 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb7 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_183 <= _pht_0_T_11;
        end else begin
          pht_0_183 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_184 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb8 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_184 <= _pht_0_T_11;
        end else begin
          pht_0_184 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_185 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hb9 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_185 <= _pht_0_T_11;
        end else begin
          pht_0_185 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_186 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hba == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_186 <= _pht_0_T_11;
        end else begin
          pht_0_186 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_187 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hbb == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_187 <= _pht_0_T_11;
        end else begin
          pht_0_187 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_188 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hbc == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_188 <= _pht_0_T_11;
        end else begin
          pht_0_188 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_189 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hbd == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_189 <= _pht_0_T_11;
        end else begin
          pht_0_189 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_190 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hbe == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_190 <= _pht_0_T_11;
        end else begin
          pht_0_190 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_191 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hbf == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_191 <= _pht_0_T_11;
        end else begin
          pht_0_191 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_192 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc0 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_192 <= _pht_0_T_11;
        end else begin
          pht_0_192 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_193 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc1 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_193 <= _pht_0_T_11;
        end else begin
          pht_0_193 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_194 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc2 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_194 <= _pht_0_T_11;
        end else begin
          pht_0_194 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_195 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc3 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_195 <= _pht_0_T_11;
        end else begin
          pht_0_195 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_196 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc4 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_196 <= _pht_0_T_11;
        end else begin
          pht_0_196 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_197 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc5 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_197 <= _pht_0_T_11;
        end else begin
          pht_0_197 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_198 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc6 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_198 <= _pht_0_T_11;
        end else begin
          pht_0_198 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_199 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc7 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_199 <= _pht_0_T_11;
        end else begin
          pht_0_199 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_200 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc8 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_200 <= _pht_0_T_11;
        end else begin
          pht_0_200 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_201 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hc9 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_201 <= _pht_0_T_11;
        end else begin
          pht_0_201 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_202 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hca == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_202 <= _pht_0_T_11;
        end else begin
          pht_0_202 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_203 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hcb == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_203 <= _pht_0_T_11;
        end else begin
          pht_0_203 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_204 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hcc == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_204 <= _pht_0_T_11;
        end else begin
          pht_0_204 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_205 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hcd == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_205 <= _pht_0_T_11;
        end else begin
          pht_0_205 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_206 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hce == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_206 <= _pht_0_T_11;
        end else begin
          pht_0_206 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_207 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hcf == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_207 <= _pht_0_T_11;
        end else begin
          pht_0_207 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_208 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd0 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_208 <= _pht_0_T_11;
        end else begin
          pht_0_208 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_209 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd1 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_209 <= _pht_0_T_11;
        end else begin
          pht_0_209 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_210 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd2 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_210 <= _pht_0_T_11;
        end else begin
          pht_0_210 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_211 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd3 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_211 <= _pht_0_T_11;
        end else begin
          pht_0_211 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_212 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd4 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_212 <= _pht_0_T_11;
        end else begin
          pht_0_212 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_213 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd5 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_213 <= _pht_0_T_11;
        end else begin
          pht_0_213 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_214 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd6 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_214 <= _pht_0_T_11;
        end else begin
          pht_0_214 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_215 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd7 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_215 <= _pht_0_T_11;
        end else begin
          pht_0_215 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_216 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd8 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_216 <= _pht_0_T_11;
        end else begin
          pht_0_216 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_217 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hd9 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_217 <= _pht_0_T_11;
        end else begin
          pht_0_217 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_218 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hda == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_218 <= _pht_0_T_11;
        end else begin
          pht_0_218 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_219 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hdb == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_219 <= _pht_0_T_11;
        end else begin
          pht_0_219 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_220 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hdc == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_220 <= _pht_0_T_11;
        end else begin
          pht_0_220 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_221 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hdd == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_221 <= _pht_0_T_11;
        end else begin
          pht_0_221 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_222 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hde == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_222 <= _pht_0_T_11;
        end else begin
          pht_0_222 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_223 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hdf == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_223 <= _pht_0_T_11;
        end else begin
          pht_0_223 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_224 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he0 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_224 <= _pht_0_T_11;
        end else begin
          pht_0_224 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_225 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he1 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_225 <= _pht_0_T_11;
        end else begin
          pht_0_225 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_226 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he2 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_226 <= _pht_0_T_11;
        end else begin
          pht_0_226 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_227 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he3 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_227 <= _pht_0_T_11;
        end else begin
          pht_0_227 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_228 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he4 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_228 <= _pht_0_T_11;
        end else begin
          pht_0_228 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_229 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he5 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_229 <= _pht_0_T_11;
        end else begin
          pht_0_229 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_230 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he6 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_230 <= _pht_0_T_11;
        end else begin
          pht_0_230 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_231 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he7 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_231 <= _pht_0_T_11;
        end else begin
          pht_0_231 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_232 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he8 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_232 <= _pht_0_T_11;
        end else begin
          pht_0_232 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_233 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'he9 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_233 <= _pht_0_T_11;
        end else begin
          pht_0_233 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_234 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hea == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_234 <= _pht_0_T_11;
        end else begin
          pht_0_234 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_235 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'heb == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_235 <= _pht_0_T_11;
        end else begin
          pht_0_235 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_236 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hec == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_236 <= _pht_0_T_11;
        end else begin
          pht_0_236 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_237 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hed == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_237 <= _pht_0_T_11;
        end else begin
          pht_0_237 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_238 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hee == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_238 <= _pht_0_T_11;
        end else begin
          pht_0_238 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_239 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hef == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_239 <= _pht_0_T_11;
        end else begin
          pht_0_239 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_240 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf0 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_240 <= _pht_0_T_11;
        end else begin
          pht_0_240 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_241 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf1 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_241 <= _pht_0_T_11;
        end else begin
          pht_0_241 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_242 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf2 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_242 <= _pht_0_T_11;
        end else begin
          pht_0_242 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_243 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf3 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_243 <= _pht_0_T_11;
        end else begin
          pht_0_243 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_244 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf4 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_244 <= _pht_0_T_11;
        end else begin
          pht_0_244 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_245 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf5 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_245 <= _pht_0_T_11;
        end else begin
          pht_0_245 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_246 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf6 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_246 <= _pht_0_T_11;
        end else begin
          pht_0_246 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_247 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf7 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_247 <= _pht_0_T_11;
        end else begin
          pht_0_247 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_248 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf8 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_248 <= _pht_0_T_11;
        end else begin
          pht_0_248 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_249 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hf9 == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_249 <= _pht_0_T_11;
        end else begin
          pht_0_249 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_250 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hfa == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_250 <= _pht_0_T_11;
        end else begin
          pht_0_250 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_251 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hfb == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_251 <= _pht_0_T_11;
        end else begin
          pht_0_251 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_252 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hfc == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_252 <= _pht_0_T_11;
        end else begin
          pht_0_252 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_253 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hfd == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_253 <= _pht_0_T_11;
        end else begin
          pht_0_253 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_254 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hfe == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_254 <= _pht_0_T_11;
        end else begin
          pht_0_254 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_0_255 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 82:25]
      if (8'hff == pht1WAddr) begin // @[bht.scala 83:25]
        if (2'h3 == _GEN_1663) begin // @[Mux.scala 81:58]
          pht_0_255 <= _pht_0_T_11;
        end else begin
          pht_0_255 <= _pht_0_T_15;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_0 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h0 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_0 <= _pht_1_T_3;
        end else begin
          pht_1_0 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_1 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h1 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_1 <= _pht_1_T_3;
        end else begin
          pht_1_1 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_2 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h2 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_2 <= _pht_1_T_3;
        end else begin
          pht_1_2 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_3 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h3 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_3 <= _pht_1_T_3;
        end else begin
          pht_1_3 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_4 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h4 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_4 <= _pht_1_T_3;
        end else begin
          pht_1_4 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_5 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h5 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_5 <= _pht_1_T_3;
        end else begin
          pht_1_5 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_6 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h6 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_6 <= _pht_1_T_3;
        end else begin
          pht_1_6 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_7 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h7 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_7 <= _pht_1_T_3;
        end else begin
          pht_1_7 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_8 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h8 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_8 <= _pht_1_T_3;
        end else begin
          pht_1_8 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_9 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h9 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_9 <= _pht_1_T_3;
        end else begin
          pht_1_9 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_10 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_10 <= _pht_1_T_3;
        end else begin
          pht_1_10 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_11 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_11 <= _pht_1_T_3;
        end else begin
          pht_1_11 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_12 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_12 <= _pht_1_T_3;
        end else begin
          pht_1_12 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_13 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_13 <= _pht_1_T_3;
        end else begin
          pht_1_13 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_14 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_14 <= _pht_1_T_3;
        end else begin
          pht_1_14 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_15 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_15 <= _pht_1_T_3;
        end else begin
          pht_1_15 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_16 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h10 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_16 <= _pht_1_T_3;
        end else begin
          pht_1_16 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_17 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h11 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_17 <= _pht_1_T_3;
        end else begin
          pht_1_17 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_18 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h12 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_18 <= _pht_1_T_3;
        end else begin
          pht_1_18 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_19 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h13 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_19 <= _pht_1_T_3;
        end else begin
          pht_1_19 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_20 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h14 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_20 <= _pht_1_T_3;
        end else begin
          pht_1_20 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_21 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h15 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_21 <= _pht_1_T_3;
        end else begin
          pht_1_21 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_22 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h16 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_22 <= _pht_1_T_3;
        end else begin
          pht_1_22 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_23 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h17 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_23 <= _pht_1_T_3;
        end else begin
          pht_1_23 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_24 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h18 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_24 <= _pht_1_T_3;
        end else begin
          pht_1_24 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_25 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h19 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_25 <= _pht_1_T_3;
        end else begin
          pht_1_25 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_26 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h1a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_26 <= _pht_1_T_3;
        end else begin
          pht_1_26 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_27 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h1b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_27 <= _pht_1_T_3;
        end else begin
          pht_1_27 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_28 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h1c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_28 <= _pht_1_T_3;
        end else begin
          pht_1_28 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_29 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h1d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_29 <= _pht_1_T_3;
        end else begin
          pht_1_29 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_30 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h1e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_30 <= _pht_1_T_3;
        end else begin
          pht_1_30 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_31 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h1f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_31 <= _pht_1_T_3;
        end else begin
          pht_1_31 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_32 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h20 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_32 <= _pht_1_T_3;
        end else begin
          pht_1_32 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_33 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h21 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_33 <= _pht_1_T_3;
        end else begin
          pht_1_33 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_34 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h22 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_34 <= _pht_1_T_3;
        end else begin
          pht_1_34 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_35 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h23 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_35 <= _pht_1_T_3;
        end else begin
          pht_1_35 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_36 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h24 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_36 <= _pht_1_T_3;
        end else begin
          pht_1_36 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_37 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h25 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_37 <= _pht_1_T_3;
        end else begin
          pht_1_37 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_38 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h26 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_38 <= _pht_1_T_3;
        end else begin
          pht_1_38 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_39 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h27 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_39 <= _pht_1_T_3;
        end else begin
          pht_1_39 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_40 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h28 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_40 <= _pht_1_T_3;
        end else begin
          pht_1_40 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_41 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h29 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_41 <= _pht_1_T_3;
        end else begin
          pht_1_41 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_42 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h2a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_42 <= _pht_1_T_3;
        end else begin
          pht_1_42 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_43 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h2b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_43 <= _pht_1_T_3;
        end else begin
          pht_1_43 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_44 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h2c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_44 <= _pht_1_T_3;
        end else begin
          pht_1_44 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_45 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h2d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_45 <= _pht_1_T_3;
        end else begin
          pht_1_45 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_46 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h2e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_46 <= _pht_1_T_3;
        end else begin
          pht_1_46 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_47 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h2f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_47 <= _pht_1_T_3;
        end else begin
          pht_1_47 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_48 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h30 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_48 <= _pht_1_T_3;
        end else begin
          pht_1_48 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_49 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h31 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_49 <= _pht_1_T_3;
        end else begin
          pht_1_49 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_50 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h32 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_50 <= _pht_1_T_3;
        end else begin
          pht_1_50 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_51 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h33 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_51 <= _pht_1_T_3;
        end else begin
          pht_1_51 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_52 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h34 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_52 <= _pht_1_T_3;
        end else begin
          pht_1_52 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_53 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h35 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_53 <= _pht_1_T_3;
        end else begin
          pht_1_53 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_54 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h36 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_54 <= _pht_1_T_3;
        end else begin
          pht_1_54 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_55 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h37 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_55 <= _pht_1_T_3;
        end else begin
          pht_1_55 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_56 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h38 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_56 <= _pht_1_T_3;
        end else begin
          pht_1_56 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_57 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h39 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_57 <= _pht_1_T_3;
        end else begin
          pht_1_57 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_58 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h3a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_58 <= _pht_1_T_3;
        end else begin
          pht_1_58 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_59 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h3b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_59 <= _pht_1_T_3;
        end else begin
          pht_1_59 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_60 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h3c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_60 <= _pht_1_T_3;
        end else begin
          pht_1_60 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_61 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h3d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_61 <= _pht_1_T_3;
        end else begin
          pht_1_61 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_62 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h3e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_62 <= _pht_1_T_3;
        end else begin
          pht_1_62 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_63 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h3f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_63 <= _pht_1_T_3;
        end else begin
          pht_1_63 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_64 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h40 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_64 <= _pht_1_T_3;
        end else begin
          pht_1_64 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_65 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h41 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_65 <= _pht_1_T_3;
        end else begin
          pht_1_65 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_66 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h42 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_66 <= _pht_1_T_3;
        end else begin
          pht_1_66 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_67 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h43 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_67 <= _pht_1_T_3;
        end else begin
          pht_1_67 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_68 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h44 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_68 <= _pht_1_T_3;
        end else begin
          pht_1_68 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_69 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h45 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_69 <= _pht_1_T_3;
        end else begin
          pht_1_69 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_70 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h46 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_70 <= _pht_1_T_3;
        end else begin
          pht_1_70 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_71 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h47 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_71 <= _pht_1_T_3;
        end else begin
          pht_1_71 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_72 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h48 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_72 <= _pht_1_T_3;
        end else begin
          pht_1_72 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_73 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h49 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_73 <= _pht_1_T_3;
        end else begin
          pht_1_73 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_74 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h4a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_74 <= _pht_1_T_3;
        end else begin
          pht_1_74 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_75 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h4b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_75 <= _pht_1_T_3;
        end else begin
          pht_1_75 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_76 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h4c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_76 <= _pht_1_T_3;
        end else begin
          pht_1_76 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_77 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h4d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_77 <= _pht_1_T_3;
        end else begin
          pht_1_77 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_78 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h4e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_78 <= _pht_1_T_3;
        end else begin
          pht_1_78 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_79 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h4f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_79 <= _pht_1_T_3;
        end else begin
          pht_1_79 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_80 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h50 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_80 <= _pht_1_T_3;
        end else begin
          pht_1_80 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_81 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h51 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_81 <= _pht_1_T_3;
        end else begin
          pht_1_81 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_82 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h52 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_82 <= _pht_1_T_3;
        end else begin
          pht_1_82 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_83 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h53 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_83 <= _pht_1_T_3;
        end else begin
          pht_1_83 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_84 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h54 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_84 <= _pht_1_T_3;
        end else begin
          pht_1_84 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_85 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h55 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_85 <= _pht_1_T_3;
        end else begin
          pht_1_85 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_86 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h56 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_86 <= _pht_1_T_3;
        end else begin
          pht_1_86 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_87 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h57 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_87 <= _pht_1_T_3;
        end else begin
          pht_1_87 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_88 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h58 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_88 <= _pht_1_T_3;
        end else begin
          pht_1_88 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_89 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h59 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_89 <= _pht_1_T_3;
        end else begin
          pht_1_89 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_90 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h5a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_90 <= _pht_1_T_3;
        end else begin
          pht_1_90 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_91 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h5b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_91 <= _pht_1_T_3;
        end else begin
          pht_1_91 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_92 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h5c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_92 <= _pht_1_T_3;
        end else begin
          pht_1_92 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_93 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h5d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_93 <= _pht_1_T_3;
        end else begin
          pht_1_93 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_94 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h5e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_94 <= _pht_1_T_3;
        end else begin
          pht_1_94 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_95 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h5f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_95 <= _pht_1_T_3;
        end else begin
          pht_1_95 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_96 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h60 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_96 <= _pht_1_T_3;
        end else begin
          pht_1_96 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_97 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h61 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_97 <= _pht_1_T_3;
        end else begin
          pht_1_97 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_98 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h62 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_98 <= _pht_1_T_3;
        end else begin
          pht_1_98 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_99 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h63 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_99 <= _pht_1_T_3;
        end else begin
          pht_1_99 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_100 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h64 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_100 <= _pht_1_T_3;
        end else begin
          pht_1_100 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_101 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h65 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_101 <= _pht_1_T_3;
        end else begin
          pht_1_101 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_102 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h66 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_102 <= _pht_1_T_3;
        end else begin
          pht_1_102 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_103 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h67 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_103 <= _pht_1_T_3;
        end else begin
          pht_1_103 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_104 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h68 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_104 <= _pht_1_T_3;
        end else begin
          pht_1_104 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_105 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h69 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_105 <= _pht_1_T_3;
        end else begin
          pht_1_105 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_106 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h6a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_106 <= _pht_1_T_3;
        end else begin
          pht_1_106 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_107 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h6b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_107 <= _pht_1_T_3;
        end else begin
          pht_1_107 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_108 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h6c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_108 <= _pht_1_T_3;
        end else begin
          pht_1_108 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_109 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h6d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_109 <= _pht_1_T_3;
        end else begin
          pht_1_109 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_110 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h6e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_110 <= _pht_1_T_3;
        end else begin
          pht_1_110 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_111 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h6f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_111 <= _pht_1_T_3;
        end else begin
          pht_1_111 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_112 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h70 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_112 <= _pht_1_T_3;
        end else begin
          pht_1_112 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_113 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h71 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_113 <= _pht_1_T_3;
        end else begin
          pht_1_113 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_114 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h72 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_114 <= _pht_1_T_3;
        end else begin
          pht_1_114 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_115 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h73 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_115 <= _pht_1_T_3;
        end else begin
          pht_1_115 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_116 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h74 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_116 <= _pht_1_T_3;
        end else begin
          pht_1_116 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_117 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h75 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_117 <= _pht_1_T_3;
        end else begin
          pht_1_117 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_118 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h76 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_118 <= _pht_1_T_3;
        end else begin
          pht_1_118 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_119 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h77 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_119 <= _pht_1_T_3;
        end else begin
          pht_1_119 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_120 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h78 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_120 <= _pht_1_T_3;
        end else begin
          pht_1_120 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_121 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h79 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_121 <= _pht_1_T_3;
        end else begin
          pht_1_121 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_122 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h7a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_122 <= _pht_1_T_3;
        end else begin
          pht_1_122 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_123 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h7b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_123 <= _pht_1_T_3;
        end else begin
          pht_1_123 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_124 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h7c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_124 <= _pht_1_T_3;
        end else begin
          pht_1_124 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_125 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h7d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_125 <= _pht_1_T_3;
        end else begin
          pht_1_125 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_126 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h7e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_126 <= _pht_1_T_3;
        end else begin
          pht_1_126 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_127 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h7f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_127 <= _pht_1_T_3;
        end else begin
          pht_1_127 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_128 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h80 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_128 <= _pht_1_T_3;
        end else begin
          pht_1_128 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_129 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h81 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_129 <= _pht_1_T_3;
        end else begin
          pht_1_129 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_130 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h82 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_130 <= _pht_1_T_3;
        end else begin
          pht_1_130 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_131 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h83 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_131 <= _pht_1_T_3;
        end else begin
          pht_1_131 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_132 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h84 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_132 <= _pht_1_T_3;
        end else begin
          pht_1_132 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_133 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h85 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_133 <= _pht_1_T_3;
        end else begin
          pht_1_133 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_134 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h86 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_134 <= _pht_1_T_3;
        end else begin
          pht_1_134 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_135 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h87 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_135 <= _pht_1_T_3;
        end else begin
          pht_1_135 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_136 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h88 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_136 <= _pht_1_T_3;
        end else begin
          pht_1_136 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_137 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h89 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_137 <= _pht_1_T_3;
        end else begin
          pht_1_137 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_138 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h8a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_138 <= _pht_1_T_3;
        end else begin
          pht_1_138 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_139 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h8b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_139 <= _pht_1_T_3;
        end else begin
          pht_1_139 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_140 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h8c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_140 <= _pht_1_T_3;
        end else begin
          pht_1_140 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_141 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h8d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_141 <= _pht_1_T_3;
        end else begin
          pht_1_141 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_142 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h8e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_142 <= _pht_1_T_3;
        end else begin
          pht_1_142 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_143 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h8f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_143 <= _pht_1_T_3;
        end else begin
          pht_1_143 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_144 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h90 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_144 <= _pht_1_T_3;
        end else begin
          pht_1_144 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_145 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h91 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_145 <= _pht_1_T_3;
        end else begin
          pht_1_145 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_146 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h92 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_146 <= _pht_1_T_3;
        end else begin
          pht_1_146 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_147 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h93 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_147 <= _pht_1_T_3;
        end else begin
          pht_1_147 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_148 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h94 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_148 <= _pht_1_T_3;
        end else begin
          pht_1_148 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_149 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h95 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_149 <= _pht_1_T_3;
        end else begin
          pht_1_149 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_150 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h96 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_150 <= _pht_1_T_3;
        end else begin
          pht_1_150 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_151 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h97 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_151 <= _pht_1_T_3;
        end else begin
          pht_1_151 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_152 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h98 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_152 <= _pht_1_T_3;
        end else begin
          pht_1_152 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_153 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h99 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_153 <= _pht_1_T_3;
        end else begin
          pht_1_153 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_154 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h9a == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_154 <= _pht_1_T_3;
        end else begin
          pht_1_154 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_155 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h9b == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_155 <= _pht_1_T_3;
        end else begin
          pht_1_155 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_156 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h9c == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_156 <= _pht_1_T_3;
        end else begin
          pht_1_156 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_157 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h9d == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_157 <= _pht_1_T_3;
        end else begin
          pht_1_157 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_158 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h9e == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_158 <= _pht_1_T_3;
        end else begin
          pht_1_158 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_159 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'h9f == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_159 <= _pht_1_T_3;
        end else begin
          pht_1_159 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_160 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha0 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_160 <= _pht_1_T_3;
        end else begin
          pht_1_160 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_161 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha1 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_161 <= _pht_1_T_3;
        end else begin
          pht_1_161 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_162 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha2 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_162 <= _pht_1_T_3;
        end else begin
          pht_1_162 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_163 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha3 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_163 <= _pht_1_T_3;
        end else begin
          pht_1_163 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_164 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha4 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_164 <= _pht_1_T_3;
        end else begin
          pht_1_164 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_165 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha5 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_165 <= _pht_1_T_3;
        end else begin
          pht_1_165 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_166 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha6 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_166 <= _pht_1_T_3;
        end else begin
          pht_1_166 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_167 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha7 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_167 <= _pht_1_T_3;
        end else begin
          pht_1_167 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_168 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha8 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_168 <= _pht_1_T_3;
        end else begin
          pht_1_168 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_169 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'ha9 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_169 <= _pht_1_T_3;
        end else begin
          pht_1_169 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_170 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'haa == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_170 <= _pht_1_T_3;
        end else begin
          pht_1_170 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_171 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hab == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_171 <= _pht_1_T_3;
        end else begin
          pht_1_171 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_172 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hac == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_172 <= _pht_1_T_3;
        end else begin
          pht_1_172 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_173 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'had == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_173 <= _pht_1_T_3;
        end else begin
          pht_1_173 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_174 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hae == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_174 <= _pht_1_T_3;
        end else begin
          pht_1_174 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_175 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'haf == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_175 <= _pht_1_T_3;
        end else begin
          pht_1_175 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_176 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb0 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_176 <= _pht_1_T_3;
        end else begin
          pht_1_176 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_177 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb1 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_177 <= _pht_1_T_3;
        end else begin
          pht_1_177 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_178 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb2 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_178 <= _pht_1_T_3;
        end else begin
          pht_1_178 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_179 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb3 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_179 <= _pht_1_T_3;
        end else begin
          pht_1_179 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_180 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb4 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_180 <= _pht_1_T_3;
        end else begin
          pht_1_180 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_181 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb5 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_181 <= _pht_1_T_3;
        end else begin
          pht_1_181 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_182 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb6 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_182 <= _pht_1_T_3;
        end else begin
          pht_1_182 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_183 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb7 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_183 <= _pht_1_T_3;
        end else begin
          pht_1_183 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_184 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb8 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_184 <= _pht_1_T_3;
        end else begin
          pht_1_184 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_185 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hb9 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_185 <= _pht_1_T_3;
        end else begin
          pht_1_185 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_186 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hba == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_186 <= _pht_1_T_3;
        end else begin
          pht_1_186 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_187 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hbb == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_187 <= _pht_1_T_3;
        end else begin
          pht_1_187 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_188 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hbc == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_188 <= _pht_1_T_3;
        end else begin
          pht_1_188 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_189 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hbd == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_189 <= _pht_1_T_3;
        end else begin
          pht_1_189 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_190 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hbe == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_190 <= _pht_1_T_3;
        end else begin
          pht_1_190 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_191 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hbf == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_191 <= _pht_1_T_3;
        end else begin
          pht_1_191 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_192 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc0 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_192 <= _pht_1_T_3;
        end else begin
          pht_1_192 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_193 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc1 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_193 <= _pht_1_T_3;
        end else begin
          pht_1_193 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_194 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc2 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_194 <= _pht_1_T_3;
        end else begin
          pht_1_194 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_195 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc3 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_195 <= _pht_1_T_3;
        end else begin
          pht_1_195 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_196 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc4 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_196 <= _pht_1_T_3;
        end else begin
          pht_1_196 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_197 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc5 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_197 <= _pht_1_T_3;
        end else begin
          pht_1_197 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_198 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc6 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_198 <= _pht_1_T_3;
        end else begin
          pht_1_198 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_199 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc7 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_199 <= _pht_1_T_3;
        end else begin
          pht_1_199 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_200 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc8 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_200 <= _pht_1_T_3;
        end else begin
          pht_1_200 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_201 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hc9 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_201 <= _pht_1_T_3;
        end else begin
          pht_1_201 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_202 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hca == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_202 <= _pht_1_T_3;
        end else begin
          pht_1_202 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_203 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hcb == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_203 <= _pht_1_T_3;
        end else begin
          pht_1_203 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_204 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hcc == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_204 <= _pht_1_T_3;
        end else begin
          pht_1_204 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_205 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hcd == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_205 <= _pht_1_T_3;
        end else begin
          pht_1_205 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_206 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hce == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_206 <= _pht_1_T_3;
        end else begin
          pht_1_206 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_207 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hcf == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_207 <= _pht_1_T_3;
        end else begin
          pht_1_207 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_208 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd0 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_208 <= _pht_1_T_3;
        end else begin
          pht_1_208 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_209 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd1 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_209 <= _pht_1_T_3;
        end else begin
          pht_1_209 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_210 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd2 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_210 <= _pht_1_T_3;
        end else begin
          pht_1_210 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_211 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd3 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_211 <= _pht_1_T_3;
        end else begin
          pht_1_211 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_212 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd4 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_212 <= _pht_1_T_3;
        end else begin
          pht_1_212 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_213 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd5 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_213 <= _pht_1_T_3;
        end else begin
          pht_1_213 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_214 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd6 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_214 <= _pht_1_T_3;
        end else begin
          pht_1_214 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_215 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd7 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_215 <= _pht_1_T_3;
        end else begin
          pht_1_215 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_216 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd8 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_216 <= _pht_1_T_3;
        end else begin
          pht_1_216 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_217 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hd9 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_217 <= _pht_1_T_3;
        end else begin
          pht_1_217 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_218 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hda == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_218 <= _pht_1_T_3;
        end else begin
          pht_1_218 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_219 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hdb == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_219 <= _pht_1_T_3;
        end else begin
          pht_1_219 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_220 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hdc == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_220 <= _pht_1_T_3;
        end else begin
          pht_1_220 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_221 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hdd == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_221 <= _pht_1_T_3;
        end else begin
          pht_1_221 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_222 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hde == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_222 <= _pht_1_T_3;
        end else begin
          pht_1_222 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_223 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hdf == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_223 <= _pht_1_T_3;
        end else begin
          pht_1_223 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_224 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he0 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_224 <= _pht_1_T_3;
        end else begin
          pht_1_224 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_225 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he1 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_225 <= _pht_1_T_3;
        end else begin
          pht_1_225 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_226 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he2 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_226 <= _pht_1_T_3;
        end else begin
          pht_1_226 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_227 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he3 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_227 <= _pht_1_T_3;
        end else begin
          pht_1_227 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_228 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he4 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_228 <= _pht_1_T_3;
        end else begin
          pht_1_228 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_229 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he5 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_229 <= _pht_1_T_3;
        end else begin
          pht_1_229 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_230 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he6 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_230 <= _pht_1_T_3;
        end else begin
          pht_1_230 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_231 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he7 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_231 <= _pht_1_T_3;
        end else begin
          pht_1_231 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_232 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he8 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_232 <= _pht_1_T_3;
        end else begin
          pht_1_232 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_233 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'he9 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_233 <= _pht_1_T_3;
        end else begin
          pht_1_233 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_234 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hea == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_234 <= _pht_1_T_3;
        end else begin
          pht_1_234 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_235 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'heb == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_235 <= _pht_1_T_3;
        end else begin
          pht_1_235 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_236 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hec == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_236 <= _pht_1_T_3;
        end else begin
          pht_1_236 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_237 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hed == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_237 <= _pht_1_T_3;
        end else begin
          pht_1_237 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_238 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hee == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_238 <= _pht_1_T_3;
        end else begin
          pht_1_238 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_239 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hef == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_239 <= _pht_1_T_3;
        end else begin
          pht_1_239 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_240 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf0 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_240 <= _pht_1_T_3;
        end else begin
          pht_1_240 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_241 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf1 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_241 <= _pht_1_T_3;
        end else begin
          pht_1_241 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_242 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf2 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_242 <= _pht_1_T_3;
        end else begin
          pht_1_242 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_243 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf3 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_243 <= _pht_1_T_3;
        end else begin
          pht_1_243 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_244 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf4 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_244 <= _pht_1_T_3;
        end else begin
          pht_1_244 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_245 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf5 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_245 <= _pht_1_T_3;
        end else begin
          pht_1_245 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_246 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf6 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_246 <= _pht_1_T_3;
        end else begin
          pht_1_246 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_247 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf7 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_247 <= _pht_1_T_3;
        end else begin
          pht_1_247 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_248 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf8 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_248 <= _pht_1_T_3;
        end else begin
          pht_1_248 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_249 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hf9 == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_249 <= _pht_1_T_3;
        end else begin
          pht_1_249 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_250 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hfa == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_250 <= _pht_1_T_3;
        end else begin
          pht_1_250 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_251 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hfb == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_251 <= _pht_1_T_3;
        end else begin
          pht_1_251 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_252 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hfc == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_252 <= _pht_1_T_3;
        end else begin
          pht_1_252 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_253 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hfd == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_253 <= _pht_1_T_3;
        end else begin
          pht_1_253 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_254 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hfe == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_254 <= _pht_1_T_3;
        end else begin
          pht_1_254 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_1_255 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 92:25]
      if (8'hff == pht1WAddr) begin // @[bht.scala 93:25]
        if (2'h3 == _GEN_1151) begin // @[Mux.scala 81:58]
          pht_1_255 <= _pht_1_T_3;
        end else begin
          pht_1_255 <= _pht_1_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_0 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h0 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_0 <= _pht_1_T_3;
        end else begin
          pht_2_0 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_1 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h1 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_1 <= _pht_1_T_3;
        end else begin
          pht_2_1 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_2 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h2 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_2 <= _pht_1_T_3;
        end else begin
          pht_2_2 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_3 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h3 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_3 <= _pht_1_T_3;
        end else begin
          pht_2_3 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_4 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h4 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_4 <= _pht_1_T_3;
        end else begin
          pht_2_4 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_5 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h5 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_5 <= _pht_1_T_3;
        end else begin
          pht_2_5 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_6 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h6 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_6 <= _pht_1_T_3;
        end else begin
          pht_2_6 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_7 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h7 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_7 <= _pht_1_T_3;
        end else begin
          pht_2_7 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_8 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h8 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_8 <= _pht_1_T_3;
        end else begin
          pht_2_8 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_9 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h9 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_9 <= _pht_1_T_3;
        end else begin
          pht_2_9 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_10 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_10 <= _pht_1_T_3;
        end else begin
          pht_2_10 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_11 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_11 <= _pht_1_T_3;
        end else begin
          pht_2_11 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_12 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_12 <= _pht_1_T_3;
        end else begin
          pht_2_12 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_13 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_13 <= _pht_1_T_3;
        end else begin
          pht_2_13 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_14 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_14 <= _pht_1_T_3;
        end else begin
          pht_2_14 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_15 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_15 <= _pht_1_T_3;
        end else begin
          pht_2_15 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_16 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h10 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_16 <= _pht_1_T_3;
        end else begin
          pht_2_16 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_17 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h11 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_17 <= _pht_1_T_3;
        end else begin
          pht_2_17 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_18 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h12 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_18 <= _pht_1_T_3;
        end else begin
          pht_2_18 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_19 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h13 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_19 <= _pht_1_T_3;
        end else begin
          pht_2_19 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_20 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h14 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_20 <= _pht_1_T_3;
        end else begin
          pht_2_20 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_21 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h15 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_21 <= _pht_1_T_3;
        end else begin
          pht_2_21 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_22 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h16 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_22 <= _pht_1_T_3;
        end else begin
          pht_2_22 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_23 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h17 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_23 <= _pht_1_T_3;
        end else begin
          pht_2_23 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_24 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h18 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_24 <= _pht_1_T_3;
        end else begin
          pht_2_24 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_25 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h19 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_25 <= _pht_1_T_3;
        end else begin
          pht_2_25 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_26 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h1a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_26 <= _pht_1_T_3;
        end else begin
          pht_2_26 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_27 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h1b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_27 <= _pht_1_T_3;
        end else begin
          pht_2_27 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_28 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h1c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_28 <= _pht_1_T_3;
        end else begin
          pht_2_28 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_29 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h1d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_29 <= _pht_1_T_3;
        end else begin
          pht_2_29 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_30 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h1e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_30 <= _pht_1_T_3;
        end else begin
          pht_2_30 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_31 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h1f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_31 <= _pht_1_T_3;
        end else begin
          pht_2_31 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_32 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h20 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_32 <= _pht_1_T_3;
        end else begin
          pht_2_32 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_33 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h21 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_33 <= _pht_1_T_3;
        end else begin
          pht_2_33 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_34 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h22 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_34 <= _pht_1_T_3;
        end else begin
          pht_2_34 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_35 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h23 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_35 <= _pht_1_T_3;
        end else begin
          pht_2_35 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_36 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h24 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_36 <= _pht_1_T_3;
        end else begin
          pht_2_36 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_37 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h25 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_37 <= _pht_1_T_3;
        end else begin
          pht_2_37 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_38 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h26 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_38 <= _pht_1_T_3;
        end else begin
          pht_2_38 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_39 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h27 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_39 <= _pht_1_T_3;
        end else begin
          pht_2_39 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_40 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h28 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_40 <= _pht_1_T_3;
        end else begin
          pht_2_40 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_41 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h29 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_41 <= _pht_1_T_3;
        end else begin
          pht_2_41 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_42 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h2a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_42 <= _pht_1_T_3;
        end else begin
          pht_2_42 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_43 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h2b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_43 <= _pht_1_T_3;
        end else begin
          pht_2_43 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_44 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h2c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_44 <= _pht_1_T_3;
        end else begin
          pht_2_44 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_45 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h2d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_45 <= _pht_1_T_3;
        end else begin
          pht_2_45 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_46 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h2e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_46 <= _pht_1_T_3;
        end else begin
          pht_2_46 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_47 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h2f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_47 <= _pht_1_T_3;
        end else begin
          pht_2_47 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_48 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h30 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_48 <= _pht_1_T_3;
        end else begin
          pht_2_48 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_49 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h31 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_49 <= _pht_1_T_3;
        end else begin
          pht_2_49 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_50 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h32 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_50 <= _pht_1_T_3;
        end else begin
          pht_2_50 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_51 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h33 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_51 <= _pht_1_T_3;
        end else begin
          pht_2_51 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_52 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h34 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_52 <= _pht_1_T_3;
        end else begin
          pht_2_52 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_53 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h35 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_53 <= _pht_1_T_3;
        end else begin
          pht_2_53 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_54 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h36 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_54 <= _pht_1_T_3;
        end else begin
          pht_2_54 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_55 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h37 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_55 <= _pht_1_T_3;
        end else begin
          pht_2_55 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_56 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h38 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_56 <= _pht_1_T_3;
        end else begin
          pht_2_56 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_57 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h39 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_57 <= _pht_1_T_3;
        end else begin
          pht_2_57 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_58 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h3a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_58 <= _pht_1_T_3;
        end else begin
          pht_2_58 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_59 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h3b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_59 <= _pht_1_T_3;
        end else begin
          pht_2_59 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_60 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h3c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_60 <= _pht_1_T_3;
        end else begin
          pht_2_60 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_61 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h3d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_61 <= _pht_1_T_3;
        end else begin
          pht_2_61 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_62 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h3e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_62 <= _pht_1_T_3;
        end else begin
          pht_2_62 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_63 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h3f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_63 <= _pht_1_T_3;
        end else begin
          pht_2_63 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_64 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h40 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_64 <= _pht_1_T_3;
        end else begin
          pht_2_64 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_65 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h41 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_65 <= _pht_1_T_3;
        end else begin
          pht_2_65 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_66 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h42 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_66 <= _pht_1_T_3;
        end else begin
          pht_2_66 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_67 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h43 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_67 <= _pht_1_T_3;
        end else begin
          pht_2_67 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_68 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h44 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_68 <= _pht_1_T_3;
        end else begin
          pht_2_68 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_69 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h45 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_69 <= _pht_1_T_3;
        end else begin
          pht_2_69 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_70 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h46 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_70 <= _pht_1_T_3;
        end else begin
          pht_2_70 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_71 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h47 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_71 <= _pht_1_T_3;
        end else begin
          pht_2_71 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_72 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h48 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_72 <= _pht_1_T_3;
        end else begin
          pht_2_72 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_73 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h49 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_73 <= _pht_1_T_3;
        end else begin
          pht_2_73 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_74 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h4a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_74 <= _pht_1_T_3;
        end else begin
          pht_2_74 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_75 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h4b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_75 <= _pht_1_T_3;
        end else begin
          pht_2_75 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_76 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h4c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_76 <= _pht_1_T_3;
        end else begin
          pht_2_76 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_77 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h4d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_77 <= _pht_1_T_3;
        end else begin
          pht_2_77 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_78 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h4e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_78 <= _pht_1_T_3;
        end else begin
          pht_2_78 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_79 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h4f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_79 <= _pht_1_T_3;
        end else begin
          pht_2_79 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_80 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h50 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_80 <= _pht_1_T_3;
        end else begin
          pht_2_80 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_81 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h51 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_81 <= _pht_1_T_3;
        end else begin
          pht_2_81 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_82 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h52 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_82 <= _pht_1_T_3;
        end else begin
          pht_2_82 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_83 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h53 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_83 <= _pht_1_T_3;
        end else begin
          pht_2_83 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_84 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h54 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_84 <= _pht_1_T_3;
        end else begin
          pht_2_84 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_85 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h55 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_85 <= _pht_1_T_3;
        end else begin
          pht_2_85 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_86 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h56 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_86 <= _pht_1_T_3;
        end else begin
          pht_2_86 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_87 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h57 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_87 <= _pht_1_T_3;
        end else begin
          pht_2_87 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_88 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h58 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_88 <= _pht_1_T_3;
        end else begin
          pht_2_88 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_89 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h59 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_89 <= _pht_1_T_3;
        end else begin
          pht_2_89 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_90 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h5a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_90 <= _pht_1_T_3;
        end else begin
          pht_2_90 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_91 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h5b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_91 <= _pht_1_T_3;
        end else begin
          pht_2_91 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_92 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h5c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_92 <= _pht_1_T_3;
        end else begin
          pht_2_92 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_93 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h5d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_93 <= _pht_1_T_3;
        end else begin
          pht_2_93 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_94 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h5e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_94 <= _pht_1_T_3;
        end else begin
          pht_2_94 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_95 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h5f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_95 <= _pht_1_T_3;
        end else begin
          pht_2_95 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_96 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h60 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_96 <= _pht_1_T_3;
        end else begin
          pht_2_96 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_97 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h61 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_97 <= _pht_1_T_3;
        end else begin
          pht_2_97 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_98 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h62 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_98 <= _pht_1_T_3;
        end else begin
          pht_2_98 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_99 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h63 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_99 <= _pht_1_T_3;
        end else begin
          pht_2_99 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_100 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h64 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_100 <= _pht_1_T_3;
        end else begin
          pht_2_100 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_101 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h65 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_101 <= _pht_1_T_3;
        end else begin
          pht_2_101 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_102 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h66 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_102 <= _pht_1_T_3;
        end else begin
          pht_2_102 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_103 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h67 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_103 <= _pht_1_T_3;
        end else begin
          pht_2_103 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_104 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h68 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_104 <= _pht_1_T_3;
        end else begin
          pht_2_104 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_105 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h69 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_105 <= _pht_1_T_3;
        end else begin
          pht_2_105 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_106 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h6a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_106 <= _pht_1_T_3;
        end else begin
          pht_2_106 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_107 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h6b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_107 <= _pht_1_T_3;
        end else begin
          pht_2_107 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_108 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h6c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_108 <= _pht_1_T_3;
        end else begin
          pht_2_108 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_109 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h6d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_109 <= _pht_1_T_3;
        end else begin
          pht_2_109 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_110 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h6e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_110 <= _pht_1_T_3;
        end else begin
          pht_2_110 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_111 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h6f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_111 <= _pht_1_T_3;
        end else begin
          pht_2_111 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_112 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h70 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_112 <= _pht_1_T_3;
        end else begin
          pht_2_112 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_113 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h71 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_113 <= _pht_1_T_3;
        end else begin
          pht_2_113 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_114 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h72 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_114 <= _pht_1_T_3;
        end else begin
          pht_2_114 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_115 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h73 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_115 <= _pht_1_T_3;
        end else begin
          pht_2_115 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_116 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h74 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_116 <= _pht_1_T_3;
        end else begin
          pht_2_116 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_117 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h75 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_117 <= _pht_1_T_3;
        end else begin
          pht_2_117 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_118 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h76 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_118 <= _pht_1_T_3;
        end else begin
          pht_2_118 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_119 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h77 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_119 <= _pht_1_T_3;
        end else begin
          pht_2_119 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_120 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h78 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_120 <= _pht_1_T_3;
        end else begin
          pht_2_120 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_121 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h79 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_121 <= _pht_1_T_3;
        end else begin
          pht_2_121 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_122 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h7a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_122 <= _pht_1_T_3;
        end else begin
          pht_2_122 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_123 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h7b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_123 <= _pht_1_T_3;
        end else begin
          pht_2_123 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_124 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h7c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_124 <= _pht_1_T_3;
        end else begin
          pht_2_124 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_125 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h7d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_125 <= _pht_1_T_3;
        end else begin
          pht_2_125 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_126 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h7e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_126 <= _pht_1_T_3;
        end else begin
          pht_2_126 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_127 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h7f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_127 <= _pht_1_T_3;
        end else begin
          pht_2_127 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_128 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h80 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_128 <= _pht_1_T_3;
        end else begin
          pht_2_128 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_129 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h81 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_129 <= _pht_1_T_3;
        end else begin
          pht_2_129 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_130 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h82 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_130 <= _pht_1_T_3;
        end else begin
          pht_2_130 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_131 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h83 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_131 <= _pht_1_T_3;
        end else begin
          pht_2_131 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_132 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h84 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_132 <= _pht_1_T_3;
        end else begin
          pht_2_132 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_133 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h85 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_133 <= _pht_1_T_3;
        end else begin
          pht_2_133 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_134 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h86 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_134 <= _pht_1_T_3;
        end else begin
          pht_2_134 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_135 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h87 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_135 <= _pht_1_T_3;
        end else begin
          pht_2_135 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_136 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h88 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_136 <= _pht_1_T_3;
        end else begin
          pht_2_136 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_137 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h89 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_137 <= _pht_1_T_3;
        end else begin
          pht_2_137 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_138 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h8a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_138 <= _pht_1_T_3;
        end else begin
          pht_2_138 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_139 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h8b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_139 <= _pht_1_T_3;
        end else begin
          pht_2_139 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_140 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h8c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_140 <= _pht_1_T_3;
        end else begin
          pht_2_140 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_141 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h8d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_141 <= _pht_1_T_3;
        end else begin
          pht_2_141 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_142 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h8e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_142 <= _pht_1_T_3;
        end else begin
          pht_2_142 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_143 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h8f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_143 <= _pht_1_T_3;
        end else begin
          pht_2_143 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_144 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h90 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_144 <= _pht_1_T_3;
        end else begin
          pht_2_144 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_145 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h91 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_145 <= _pht_1_T_3;
        end else begin
          pht_2_145 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_146 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h92 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_146 <= _pht_1_T_3;
        end else begin
          pht_2_146 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_147 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h93 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_147 <= _pht_1_T_3;
        end else begin
          pht_2_147 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_148 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h94 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_148 <= _pht_1_T_3;
        end else begin
          pht_2_148 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_149 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h95 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_149 <= _pht_1_T_3;
        end else begin
          pht_2_149 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_150 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h96 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_150 <= _pht_1_T_3;
        end else begin
          pht_2_150 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_151 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h97 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_151 <= _pht_1_T_3;
        end else begin
          pht_2_151 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_152 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h98 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_152 <= _pht_1_T_3;
        end else begin
          pht_2_152 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_153 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h99 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_153 <= _pht_1_T_3;
        end else begin
          pht_2_153 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_154 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h9a == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_154 <= _pht_1_T_3;
        end else begin
          pht_2_154 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_155 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h9b == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_155 <= _pht_1_T_3;
        end else begin
          pht_2_155 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_156 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h9c == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_156 <= _pht_1_T_3;
        end else begin
          pht_2_156 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_157 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h9d == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_157 <= _pht_1_T_3;
        end else begin
          pht_2_157 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_158 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h9e == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_158 <= _pht_1_T_3;
        end else begin
          pht_2_158 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_159 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'h9f == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_159 <= _pht_1_T_3;
        end else begin
          pht_2_159 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_160 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha0 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_160 <= _pht_1_T_3;
        end else begin
          pht_2_160 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_161 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha1 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_161 <= _pht_1_T_3;
        end else begin
          pht_2_161 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_162 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha2 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_162 <= _pht_1_T_3;
        end else begin
          pht_2_162 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_163 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha3 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_163 <= _pht_1_T_3;
        end else begin
          pht_2_163 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_164 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha4 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_164 <= _pht_1_T_3;
        end else begin
          pht_2_164 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_165 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha5 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_165 <= _pht_1_T_3;
        end else begin
          pht_2_165 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_166 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha6 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_166 <= _pht_1_T_3;
        end else begin
          pht_2_166 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_167 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha7 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_167 <= _pht_1_T_3;
        end else begin
          pht_2_167 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_168 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha8 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_168 <= _pht_1_T_3;
        end else begin
          pht_2_168 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_169 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'ha9 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_169 <= _pht_1_T_3;
        end else begin
          pht_2_169 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_170 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'haa == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_170 <= _pht_1_T_3;
        end else begin
          pht_2_170 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_171 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hab == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_171 <= _pht_1_T_3;
        end else begin
          pht_2_171 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_172 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hac == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_172 <= _pht_1_T_3;
        end else begin
          pht_2_172 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_173 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'had == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_173 <= _pht_1_T_3;
        end else begin
          pht_2_173 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_174 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hae == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_174 <= _pht_1_T_3;
        end else begin
          pht_2_174 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_175 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'haf == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_175 <= _pht_1_T_3;
        end else begin
          pht_2_175 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_176 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb0 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_176 <= _pht_1_T_3;
        end else begin
          pht_2_176 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_177 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb1 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_177 <= _pht_1_T_3;
        end else begin
          pht_2_177 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_178 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb2 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_178 <= _pht_1_T_3;
        end else begin
          pht_2_178 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_179 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb3 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_179 <= _pht_1_T_3;
        end else begin
          pht_2_179 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_180 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb4 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_180 <= _pht_1_T_3;
        end else begin
          pht_2_180 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_181 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb5 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_181 <= _pht_1_T_3;
        end else begin
          pht_2_181 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_182 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb6 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_182 <= _pht_1_T_3;
        end else begin
          pht_2_182 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_183 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb7 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_183 <= _pht_1_T_3;
        end else begin
          pht_2_183 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_184 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb8 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_184 <= _pht_1_T_3;
        end else begin
          pht_2_184 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_185 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hb9 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_185 <= _pht_1_T_3;
        end else begin
          pht_2_185 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_186 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hba == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_186 <= _pht_1_T_3;
        end else begin
          pht_2_186 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_187 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hbb == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_187 <= _pht_1_T_3;
        end else begin
          pht_2_187 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_188 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hbc == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_188 <= _pht_1_T_3;
        end else begin
          pht_2_188 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_189 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hbd == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_189 <= _pht_1_T_3;
        end else begin
          pht_2_189 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_190 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hbe == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_190 <= _pht_1_T_3;
        end else begin
          pht_2_190 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_191 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hbf == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_191 <= _pht_1_T_3;
        end else begin
          pht_2_191 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_192 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc0 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_192 <= _pht_1_T_3;
        end else begin
          pht_2_192 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_193 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc1 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_193 <= _pht_1_T_3;
        end else begin
          pht_2_193 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_194 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc2 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_194 <= _pht_1_T_3;
        end else begin
          pht_2_194 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_195 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc3 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_195 <= _pht_1_T_3;
        end else begin
          pht_2_195 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_196 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc4 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_196 <= _pht_1_T_3;
        end else begin
          pht_2_196 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_197 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc5 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_197 <= _pht_1_T_3;
        end else begin
          pht_2_197 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_198 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc6 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_198 <= _pht_1_T_3;
        end else begin
          pht_2_198 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_199 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc7 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_199 <= _pht_1_T_3;
        end else begin
          pht_2_199 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_200 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc8 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_200 <= _pht_1_T_3;
        end else begin
          pht_2_200 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_201 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hc9 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_201 <= _pht_1_T_3;
        end else begin
          pht_2_201 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_202 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hca == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_202 <= _pht_1_T_3;
        end else begin
          pht_2_202 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_203 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hcb == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_203 <= _pht_1_T_3;
        end else begin
          pht_2_203 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_204 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hcc == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_204 <= _pht_1_T_3;
        end else begin
          pht_2_204 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_205 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hcd == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_205 <= _pht_1_T_3;
        end else begin
          pht_2_205 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_206 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hce == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_206 <= _pht_1_T_3;
        end else begin
          pht_2_206 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_207 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hcf == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_207 <= _pht_1_T_3;
        end else begin
          pht_2_207 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_208 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd0 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_208 <= _pht_1_T_3;
        end else begin
          pht_2_208 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_209 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd1 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_209 <= _pht_1_T_3;
        end else begin
          pht_2_209 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_210 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd2 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_210 <= _pht_1_T_3;
        end else begin
          pht_2_210 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_211 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd3 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_211 <= _pht_1_T_3;
        end else begin
          pht_2_211 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_212 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd4 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_212 <= _pht_1_T_3;
        end else begin
          pht_2_212 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_213 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd5 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_213 <= _pht_1_T_3;
        end else begin
          pht_2_213 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_214 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd6 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_214 <= _pht_1_T_3;
        end else begin
          pht_2_214 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_215 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd7 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_215 <= _pht_1_T_3;
        end else begin
          pht_2_215 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_216 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd8 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_216 <= _pht_1_T_3;
        end else begin
          pht_2_216 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_217 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hd9 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_217 <= _pht_1_T_3;
        end else begin
          pht_2_217 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_218 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hda == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_218 <= _pht_1_T_3;
        end else begin
          pht_2_218 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_219 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hdb == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_219 <= _pht_1_T_3;
        end else begin
          pht_2_219 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_220 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hdc == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_220 <= _pht_1_T_3;
        end else begin
          pht_2_220 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_221 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hdd == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_221 <= _pht_1_T_3;
        end else begin
          pht_2_221 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_222 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hde == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_222 <= _pht_1_T_3;
        end else begin
          pht_2_222 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_223 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hdf == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_223 <= _pht_1_T_3;
        end else begin
          pht_2_223 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_224 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he0 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_224 <= _pht_1_T_3;
        end else begin
          pht_2_224 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_225 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he1 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_225 <= _pht_1_T_3;
        end else begin
          pht_2_225 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_226 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he2 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_226 <= _pht_1_T_3;
        end else begin
          pht_2_226 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_227 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he3 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_227 <= _pht_1_T_3;
        end else begin
          pht_2_227 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_228 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he4 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_228 <= _pht_1_T_3;
        end else begin
          pht_2_228 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_229 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he5 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_229 <= _pht_1_T_3;
        end else begin
          pht_2_229 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_230 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he6 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_230 <= _pht_1_T_3;
        end else begin
          pht_2_230 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_231 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he7 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_231 <= _pht_1_T_3;
        end else begin
          pht_2_231 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_232 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he8 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_232 <= _pht_1_T_3;
        end else begin
          pht_2_232 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_233 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'he9 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_233 <= _pht_1_T_3;
        end else begin
          pht_2_233 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_234 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hea == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_234 <= _pht_1_T_3;
        end else begin
          pht_2_234 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_235 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'heb == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_235 <= _pht_1_T_3;
        end else begin
          pht_2_235 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_236 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hec == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_236 <= _pht_1_T_3;
        end else begin
          pht_2_236 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_237 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hed == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_237 <= _pht_1_T_3;
        end else begin
          pht_2_237 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_238 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hee == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_238 <= _pht_1_T_3;
        end else begin
          pht_2_238 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_239 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hef == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_239 <= _pht_1_T_3;
        end else begin
          pht_2_239 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_240 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf0 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_240 <= _pht_1_T_3;
        end else begin
          pht_2_240 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_241 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf1 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_241 <= _pht_1_T_3;
        end else begin
          pht_2_241 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_242 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf2 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_242 <= _pht_1_T_3;
        end else begin
          pht_2_242 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_243 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf3 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_243 <= _pht_1_T_3;
        end else begin
          pht_2_243 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_244 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf4 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_244 <= _pht_1_T_3;
        end else begin
          pht_2_244 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_245 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf5 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_245 <= _pht_1_T_3;
        end else begin
          pht_2_245 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_246 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf6 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_246 <= _pht_1_T_3;
        end else begin
          pht_2_246 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_247 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf7 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_247 <= _pht_1_T_3;
        end else begin
          pht_2_247 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_248 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf8 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_248 <= _pht_1_T_3;
        end else begin
          pht_2_248 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_249 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hf9 == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_249 <= _pht_1_T_3;
        end else begin
          pht_2_249 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_250 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hfa == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_250 <= _pht_1_T_3;
        end else begin
          pht_2_250 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_251 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hfb == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_251 <= _pht_1_T_3;
        end else begin
          pht_2_251 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_252 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hfc == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_252 <= _pht_1_T_3;
        end else begin
          pht_2_252 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_253 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hfd == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_253 <= _pht_1_T_3;
        end else begin
          pht_2_253 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_254 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hfe == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_254 <= _pht_1_T_3;
        end else begin
          pht_2_254 <= _pht_2_T_7;
        end
      end
    end
    if (reset) begin // @[bht.scala 53:22]
      pht_2_255 <= 2'h1; // @[bht.scala 53:22]
    end else if (io_takenValid) begin // @[bht.scala 100:25]
      if (8'hff == pht2WAddr) begin // @[bht.scala 101:25]
        if (2'h3 == _GEN_1407) begin // @[Mux.scala 81:58]
          pht_2_255 <= _pht_1_T_3;
        end else begin
          pht_2_255 <= _pht_2_T_7;
        end
      end
    end
    io_ready_REG <= io_valid; // @[bht.scala 64:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ghr = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  bht_0 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  bht_1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  bht_2 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  bht_3 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  bht_4 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  bht_5 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  bht_6 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  bht_7 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  bht_8 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  bht_9 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  bht_10 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  bht_11 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  bht_12 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  bht_13 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  bht_14 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  bht_15 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  bht_16 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  bht_17 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  bht_18 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  bht_19 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  bht_20 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  bht_21 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  bht_22 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  bht_23 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  bht_24 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  bht_25 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  bht_26 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  bht_27 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  bht_28 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  bht_29 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  bht_30 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  bht_31 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  bht_32 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  bht_33 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  bht_34 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  bht_35 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  bht_36 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  bht_37 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  bht_38 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  bht_39 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  bht_40 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  bht_41 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  bht_42 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  bht_43 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  bht_44 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  bht_45 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  bht_46 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  bht_47 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  bht_48 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  bht_49 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  bht_50 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  bht_51 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  bht_52 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  bht_53 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  bht_54 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  bht_55 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  bht_56 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  bht_57 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  bht_58 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  bht_59 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  bht_60 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  bht_61 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  bht_62 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  bht_63 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  pht_0_0 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pht_0_1 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pht_0_2 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pht_0_3 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pht_0_4 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pht_0_5 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pht_0_6 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pht_0_7 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pht_0_8 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pht_0_9 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pht_0_10 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pht_0_11 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pht_0_12 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pht_0_13 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pht_0_14 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  pht_0_15 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  pht_0_16 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  pht_0_17 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  pht_0_18 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  pht_0_19 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  pht_0_20 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  pht_0_21 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  pht_0_22 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  pht_0_23 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  pht_0_24 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  pht_0_25 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  pht_0_26 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  pht_0_27 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  pht_0_28 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  pht_0_29 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  pht_0_30 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  pht_0_31 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  pht_0_32 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  pht_0_33 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  pht_0_34 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  pht_0_35 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  pht_0_36 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  pht_0_37 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  pht_0_38 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  pht_0_39 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  pht_0_40 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  pht_0_41 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  pht_0_42 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  pht_0_43 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  pht_0_44 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  pht_0_45 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  pht_0_46 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  pht_0_47 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  pht_0_48 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  pht_0_49 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  pht_0_50 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  pht_0_51 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  pht_0_52 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  pht_0_53 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  pht_0_54 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  pht_0_55 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  pht_0_56 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  pht_0_57 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  pht_0_58 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  pht_0_59 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  pht_0_60 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  pht_0_61 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  pht_0_62 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  pht_0_63 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  pht_0_64 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  pht_0_65 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  pht_0_66 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  pht_0_67 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  pht_0_68 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  pht_0_69 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  pht_0_70 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  pht_0_71 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  pht_0_72 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  pht_0_73 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  pht_0_74 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  pht_0_75 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  pht_0_76 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  pht_0_77 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  pht_0_78 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  pht_0_79 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  pht_0_80 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  pht_0_81 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  pht_0_82 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  pht_0_83 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  pht_0_84 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  pht_0_85 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  pht_0_86 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  pht_0_87 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  pht_0_88 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  pht_0_89 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  pht_0_90 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  pht_0_91 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  pht_0_92 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  pht_0_93 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  pht_0_94 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  pht_0_95 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  pht_0_96 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  pht_0_97 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  pht_0_98 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  pht_0_99 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  pht_0_100 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  pht_0_101 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  pht_0_102 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  pht_0_103 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  pht_0_104 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  pht_0_105 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  pht_0_106 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  pht_0_107 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  pht_0_108 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  pht_0_109 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  pht_0_110 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  pht_0_111 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  pht_0_112 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  pht_0_113 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  pht_0_114 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  pht_0_115 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  pht_0_116 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  pht_0_117 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  pht_0_118 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  pht_0_119 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  pht_0_120 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  pht_0_121 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  pht_0_122 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  pht_0_123 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  pht_0_124 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  pht_0_125 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  pht_0_126 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  pht_0_127 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  pht_0_128 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  pht_0_129 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  pht_0_130 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  pht_0_131 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  pht_0_132 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  pht_0_133 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  pht_0_134 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  pht_0_135 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  pht_0_136 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  pht_0_137 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  pht_0_138 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  pht_0_139 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  pht_0_140 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  pht_0_141 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  pht_0_142 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  pht_0_143 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  pht_0_144 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  pht_0_145 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  pht_0_146 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  pht_0_147 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  pht_0_148 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  pht_0_149 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  pht_0_150 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  pht_0_151 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  pht_0_152 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  pht_0_153 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  pht_0_154 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  pht_0_155 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  pht_0_156 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  pht_0_157 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  pht_0_158 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  pht_0_159 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  pht_0_160 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  pht_0_161 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  pht_0_162 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  pht_0_163 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  pht_0_164 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  pht_0_165 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  pht_0_166 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  pht_0_167 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  pht_0_168 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  pht_0_169 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  pht_0_170 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  pht_0_171 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  pht_0_172 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  pht_0_173 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  pht_0_174 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  pht_0_175 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  pht_0_176 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  pht_0_177 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  pht_0_178 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  pht_0_179 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  pht_0_180 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  pht_0_181 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  pht_0_182 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  pht_0_183 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  pht_0_184 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  pht_0_185 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  pht_0_186 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  pht_0_187 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  pht_0_188 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  pht_0_189 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  pht_0_190 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  pht_0_191 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  pht_0_192 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  pht_0_193 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  pht_0_194 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  pht_0_195 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  pht_0_196 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  pht_0_197 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  pht_0_198 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  pht_0_199 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  pht_0_200 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  pht_0_201 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  pht_0_202 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  pht_0_203 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  pht_0_204 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  pht_0_205 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  pht_0_206 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  pht_0_207 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  pht_0_208 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  pht_0_209 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  pht_0_210 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  pht_0_211 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  pht_0_212 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  pht_0_213 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  pht_0_214 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  pht_0_215 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  pht_0_216 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  pht_0_217 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  pht_0_218 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  pht_0_219 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  pht_0_220 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  pht_0_221 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  pht_0_222 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  pht_0_223 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  pht_0_224 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  pht_0_225 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  pht_0_226 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  pht_0_227 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  pht_0_228 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  pht_0_229 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  pht_0_230 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  pht_0_231 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  pht_0_232 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  pht_0_233 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  pht_0_234 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  pht_0_235 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  pht_0_236 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  pht_0_237 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  pht_0_238 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  pht_0_239 = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  pht_0_240 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  pht_0_241 = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  pht_0_242 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  pht_0_243 = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  pht_0_244 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  pht_0_245 = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  pht_0_246 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  pht_0_247 = _RAND_312[1:0];
  _RAND_313 = {1{`RANDOM}};
  pht_0_248 = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  pht_0_249 = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  pht_0_250 = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  pht_0_251 = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  pht_0_252 = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  pht_0_253 = _RAND_318[1:0];
  _RAND_319 = {1{`RANDOM}};
  pht_0_254 = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  pht_0_255 = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  pht_1_0 = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  pht_1_1 = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  pht_1_2 = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  pht_1_3 = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  pht_1_4 = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  pht_1_5 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  pht_1_6 = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  pht_1_7 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  pht_1_8 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  pht_1_9 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  pht_1_10 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  pht_1_11 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  pht_1_12 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  pht_1_13 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  pht_1_14 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  pht_1_15 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  pht_1_16 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  pht_1_17 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  pht_1_18 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  pht_1_19 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  pht_1_20 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  pht_1_21 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  pht_1_22 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  pht_1_23 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  pht_1_24 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  pht_1_25 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  pht_1_26 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  pht_1_27 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  pht_1_28 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  pht_1_29 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  pht_1_30 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  pht_1_31 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  pht_1_32 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  pht_1_33 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  pht_1_34 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  pht_1_35 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  pht_1_36 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  pht_1_37 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  pht_1_38 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  pht_1_39 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  pht_1_40 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  pht_1_41 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  pht_1_42 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  pht_1_43 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  pht_1_44 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  pht_1_45 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  pht_1_46 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  pht_1_47 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  pht_1_48 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  pht_1_49 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  pht_1_50 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  pht_1_51 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  pht_1_52 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  pht_1_53 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  pht_1_54 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  pht_1_55 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  pht_1_56 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  pht_1_57 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  pht_1_58 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  pht_1_59 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  pht_1_60 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  pht_1_61 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  pht_1_62 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  pht_1_63 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  pht_1_64 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  pht_1_65 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  pht_1_66 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  pht_1_67 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  pht_1_68 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  pht_1_69 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  pht_1_70 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  pht_1_71 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  pht_1_72 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  pht_1_73 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  pht_1_74 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  pht_1_75 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  pht_1_76 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  pht_1_77 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  pht_1_78 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  pht_1_79 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  pht_1_80 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  pht_1_81 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  pht_1_82 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  pht_1_83 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  pht_1_84 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  pht_1_85 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  pht_1_86 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  pht_1_87 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  pht_1_88 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  pht_1_89 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  pht_1_90 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  pht_1_91 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  pht_1_92 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  pht_1_93 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  pht_1_94 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  pht_1_95 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  pht_1_96 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  pht_1_97 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  pht_1_98 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  pht_1_99 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  pht_1_100 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  pht_1_101 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  pht_1_102 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  pht_1_103 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  pht_1_104 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  pht_1_105 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  pht_1_106 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  pht_1_107 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  pht_1_108 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  pht_1_109 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  pht_1_110 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  pht_1_111 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  pht_1_112 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  pht_1_113 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  pht_1_114 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  pht_1_115 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  pht_1_116 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  pht_1_117 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  pht_1_118 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  pht_1_119 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  pht_1_120 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  pht_1_121 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  pht_1_122 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  pht_1_123 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  pht_1_124 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  pht_1_125 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  pht_1_126 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  pht_1_127 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  pht_1_128 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  pht_1_129 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  pht_1_130 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  pht_1_131 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  pht_1_132 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  pht_1_133 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  pht_1_134 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  pht_1_135 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  pht_1_136 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  pht_1_137 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  pht_1_138 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  pht_1_139 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  pht_1_140 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  pht_1_141 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  pht_1_142 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  pht_1_143 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  pht_1_144 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  pht_1_145 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  pht_1_146 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  pht_1_147 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  pht_1_148 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  pht_1_149 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  pht_1_150 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  pht_1_151 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  pht_1_152 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  pht_1_153 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  pht_1_154 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  pht_1_155 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  pht_1_156 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  pht_1_157 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  pht_1_158 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  pht_1_159 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  pht_1_160 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  pht_1_161 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  pht_1_162 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  pht_1_163 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  pht_1_164 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  pht_1_165 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  pht_1_166 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  pht_1_167 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  pht_1_168 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  pht_1_169 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  pht_1_170 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  pht_1_171 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  pht_1_172 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  pht_1_173 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  pht_1_174 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  pht_1_175 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  pht_1_176 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  pht_1_177 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  pht_1_178 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  pht_1_179 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  pht_1_180 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  pht_1_181 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  pht_1_182 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  pht_1_183 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  pht_1_184 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  pht_1_185 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  pht_1_186 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  pht_1_187 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  pht_1_188 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  pht_1_189 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  pht_1_190 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  pht_1_191 = _RAND_512[1:0];
  _RAND_513 = {1{`RANDOM}};
  pht_1_192 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  pht_1_193 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  pht_1_194 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  pht_1_195 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  pht_1_196 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  pht_1_197 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  pht_1_198 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  pht_1_199 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  pht_1_200 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  pht_1_201 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  pht_1_202 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  pht_1_203 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  pht_1_204 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  pht_1_205 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  pht_1_206 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  pht_1_207 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  pht_1_208 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  pht_1_209 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  pht_1_210 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  pht_1_211 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  pht_1_212 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  pht_1_213 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  pht_1_214 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  pht_1_215 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  pht_1_216 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  pht_1_217 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  pht_1_218 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  pht_1_219 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  pht_1_220 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  pht_1_221 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  pht_1_222 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  pht_1_223 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  pht_1_224 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  pht_1_225 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  pht_1_226 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  pht_1_227 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  pht_1_228 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  pht_1_229 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  pht_1_230 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  pht_1_231 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  pht_1_232 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  pht_1_233 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  pht_1_234 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  pht_1_235 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  pht_1_236 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  pht_1_237 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  pht_1_238 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  pht_1_239 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  pht_1_240 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  pht_1_241 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  pht_1_242 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  pht_1_243 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  pht_1_244 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  pht_1_245 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  pht_1_246 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  pht_1_247 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  pht_1_248 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  pht_1_249 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  pht_1_250 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  pht_1_251 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  pht_1_252 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  pht_1_253 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  pht_1_254 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  pht_1_255 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  pht_2_0 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  pht_2_1 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  pht_2_2 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  pht_2_3 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  pht_2_4 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  pht_2_5 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  pht_2_6 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  pht_2_7 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  pht_2_8 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  pht_2_9 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  pht_2_10 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  pht_2_11 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  pht_2_12 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  pht_2_13 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  pht_2_14 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  pht_2_15 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  pht_2_16 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  pht_2_17 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  pht_2_18 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  pht_2_19 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  pht_2_20 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  pht_2_21 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  pht_2_22 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  pht_2_23 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  pht_2_24 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  pht_2_25 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  pht_2_26 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  pht_2_27 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  pht_2_28 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  pht_2_29 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  pht_2_30 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  pht_2_31 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  pht_2_32 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  pht_2_33 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  pht_2_34 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  pht_2_35 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  pht_2_36 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  pht_2_37 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  pht_2_38 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  pht_2_39 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  pht_2_40 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  pht_2_41 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  pht_2_42 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  pht_2_43 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  pht_2_44 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  pht_2_45 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  pht_2_46 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  pht_2_47 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  pht_2_48 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  pht_2_49 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  pht_2_50 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  pht_2_51 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  pht_2_52 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  pht_2_53 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  pht_2_54 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  pht_2_55 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  pht_2_56 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  pht_2_57 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  pht_2_58 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  pht_2_59 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  pht_2_60 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  pht_2_61 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  pht_2_62 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  pht_2_63 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  pht_2_64 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  pht_2_65 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  pht_2_66 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  pht_2_67 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  pht_2_68 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  pht_2_69 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  pht_2_70 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  pht_2_71 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  pht_2_72 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  pht_2_73 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  pht_2_74 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  pht_2_75 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  pht_2_76 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  pht_2_77 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  pht_2_78 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  pht_2_79 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  pht_2_80 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  pht_2_81 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  pht_2_82 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  pht_2_83 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  pht_2_84 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  pht_2_85 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  pht_2_86 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  pht_2_87 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  pht_2_88 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  pht_2_89 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  pht_2_90 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  pht_2_91 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  pht_2_92 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  pht_2_93 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  pht_2_94 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  pht_2_95 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  pht_2_96 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  pht_2_97 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  pht_2_98 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  pht_2_99 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  pht_2_100 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  pht_2_101 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  pht_2_102 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  pht_2_103 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  pht_2_104 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  pht_2_105 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  pht_2_106 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  pht_2_107 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  pht_2_108 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  pht_2_109 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  pht_2_110 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  pht_2_111 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  pht_2_112 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  pht_2_113 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  pht_2_114 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  pht_2_115 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  pht_2_116 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  pht_2_117 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  pht_2_118 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  pht_2_119 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  pht_2_120 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  pht_2_121 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  pht_2_122 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  pht_2_123 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  pht_2_124 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  pht_2_125 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  pht_2_126 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  pht_2_127 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  pht_2_128 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  pht_2_129 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  pht_2_130 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  pht_2_131 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  pht_2_132 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  pht_2_133 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  pht_2_134 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  pht_2_135 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  pht_2_136 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  pht_2_137 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  pht_2_138 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  pht_2_139 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  pht_2_140 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  pht_2_141 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  pht_2_142 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  pht_2_143 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  pht_2_144 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  pht_2_145 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  pht_2_146 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  pht_2_147 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  pht_2_148 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  pht_2_149 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  pht_2_150 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  pht_2_151 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  pht_2_152 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  pht_2_153 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  pht_2_154 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  pht_2_155 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  pht_2_156 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  pht_2_157 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  pht_2_158 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  pht_2_159 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  pht_2_160 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  pht_2_161 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  pht_2_162 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  pht_2_163 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  pht_2_164 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  pht_2_165 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  pht_2_166 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  pht_2_167 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  pht_2_168 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  pht_2_169 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  pht_2_170 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  pht_2_171 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  pht_2_172 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  pht_2_173 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  pht_2_174 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  pht_2_175 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  pht_2_176 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  pht_2_177 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  pht_2_178 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  pht_2_179 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  pht_2_180 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  pht_2_181 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  pht_2_182 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  pht_2_183 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  pht_2_184 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  pht_2_185 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  pht_2_186 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  pht_2_187 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  pht_2_188 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  pht_2_189 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  pht_2_190 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  pht_2_191 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  pht_2_192 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  pht_2_193 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  pht_2_194 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  pht_2_195 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  pht_2_196 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  pht_2_197 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  pht_2_198 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  pht_2_199 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  pht_2_200 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  pht_2_201 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  pht_2_202 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  pht_2_203 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  pht_2_204 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  pht_2_205 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  pht_2_206 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  pht_2_207 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  pht_2_208 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  pht_2_209 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  pht_2_210 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  pht_2_211 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  pht_2_212 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  pht_2_213 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  pht_2_214 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  pht_2_215 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  pht_2_216 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  pht_2_217 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  pht_2_218 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  pht_2_219 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  pht_2_220 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  pht_2_221 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  pht_2_222 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  pht_2_223 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  pht_2_224 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  pht_2_225 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  pht_2_226 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  pht_2_227 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  pht_2_228 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  pht_2_229 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  pht_2_230 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  pht_2_231 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  pht_2_232 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  pht_2_233 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  pht_2_234 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  pht_2_235 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  pht_2_236 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  pht_2_237 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  pht_2_238 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  pht_2_239 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  pht_2_240 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  pht_2_241 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  pht_2_242 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  pht_2_243 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  pht_2_244 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  pht_2_245 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  pht_2_246 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  pht_2_247 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  pht_2_248 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  pht_2_249 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  pht_2_250 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  pht_2_251 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  pht_2_252 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  pht_2_253 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  pht_2_254 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  pht_2_255 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  io_ready_REG = _RAND_833[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
